��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+�������;���ȹ�v{2� ۝ߎ#�W�ӂ����ݠ��>_g5���t͉□K2���Ec�ſ��`\_��cW��Y���NB��*�!�#-/�����0�����e	�.ZDG����g/G�lз������s�VS�]��	�_,��ܳЅ2꩙Ō��M=룯+�&HfUk�@��%��.���cm���pZ�^�&]C��l�QQ���UicM���*�qz��ZU�^u]�2�=>���J��מ�#�^Ķ���l�\*l^���F��A��N�QI�������T�xĞ��pǚ z���4��)�7�z�wcl9du�f,u���� OK���ي�H�I� ��l��.O � F�		�,& �����ͽ�`� 7�(������,\��S�!�4��ݮW���l@����1`q�f�>�U�g��E�����a�md������N���+���+���}���t�
I��-�&���I;c�C&�Q�J���5땕�?�Z|D�YP��e�|*���#܉B,��S�(����L���͙�p�&d�d�d;B�Hᨷ�ǻ��qa�+���  YEɃ��)=��������Hr߈�/G�S�>������`0&	�wu^+�#C)H�C��f�k��U�lv��v��״KOgC�Ѯx��X���8�xh��]�
�J\:�68i���Z�O	G���[s�B:�E�6M�x=	��Y�hw�946�֊0�緪&�td����q��)6�wqx��L53e�ș@h)�}Z
{�z;�L� �HW�o��>�������T��Ք�x���W��#�϶�s��B�t~��%B8��S�96C�/T��C<����!���:o��T�v�3R0`j�>��V阜��[���EU��J����dL/t��k,`��:RJ�B�I���'�9)�@j3VӘ��Jzxf���:��t�	��-(ȡ(�7���c&�"^�Y������b˓������(Xu�2'���q���N�t�#�ޜi�����'R4������(����7;��+�y���p��O薟������?�8�$�Q�o��,�c�6�PST���'�T����9gL���k?�`Zb9DTd��mL�l[����qJ�PK� �G���P#:O��̀VwG#�5b��[�69/z=�	 e,�5k@�v��J�5��q, ���8>�Ƈ�H��^*�[���u/l�Y�w`�6������Jw�:��+S�!����4�F*�X�z5<A��������ө�&W���0��`~	[Y۳��d��V���]���+@��=K����N������I�7�bV0 Z�?0�\)�����4O?d 3�!ث�7%00��K�J���wbKMB��\R�Q�FW4���^�<��[XÛx���2K.�<��_��7eTճ�X�z�U�ԂnP$R��D�(o��Aٽ��gl�ӊt�[}B���^���f� ���pc�vX��#�*�M�]��[=Bm��J��jUT�p��n��2쒏�zu�F��R�<���`=tީ�Й"��Q����J7��n�*技y��d2����@4�D9�~:���dd��v����~�cѫ�'���zL�/N^�`��V�ݎ`,JxZ^��������g)�D�?�~�e�zuw����?���J%�x�їb/{φql�H�V
	�����1,L��A�a�����R���VLU�-��]כ��v� �Ə~c��瑳_<XmVAW@�n���"��P��OK��\j�[�Pt�"���Љa9/b#?�a�V�Wv �B6����[
�wp�tg	���v�zH����"P9����$���2�޹L���-�2�tIW����o�ck�7����`5VѯM0]�^K%g����;{{�G?����R8�vQ��>���mJ�/�k�G�G�+��\@���O���o	���`>
fI�H�F"�+��{q�D�:��Pjt:�:�i������J+�,]��DQ4��sjjK(�,ӷ��$į~/>&�2�ԪL�I6;-"�S�&1�RZ�H,�*>2x`��yL��_ܺ��'i��`��������x����A~���{��ܸ]�]���v�o��Ӡj�9�CO-ETlRY�ǁ�
ك�{>%E�p�o�Oغ���`y�Ԡ���,#��i$��"�v���CNA�lk7�����t++e(fg$�ݳ��K���d�����dy�?N6�LON�o�.ur��G��cP+�P�^�Ʌ��*v�7Zs���.R�v��*:�ׁ�#j�&�v�p���	=����0l���P��������e��i�;Ǻ����?�T��+���`�!���-��-!0OXF��d�CwHS�<�hW7�oGHZR=6�8�������4�b���glDg�v�Gc��be��e�u���X�ec��f2���`A;�{�&����'��[xxݭ�ݽ1����Y�>��K7��N��;c�v \�~R�����(,c�A ϱH�����P�H]�''�������� ��TZ��d�/NG���A�ӷ��^�UX��6�e�W���� ˥����u:��3�ὼ��a.�紤ux�zU�{l��� ��	��K�2!��\��Q���K_Ö� �$����s0u��r����.y������&���!�̪����˯n6)�P�E�)��:��.�%y�#���9?f����ݡ1�_�X�Y+����1ԋH�	:�G� �Fa7����]V��o  ������6�0_��"��X�p��E-��5��~�)��!;�ȍ�������B����o���F<�)�d���;a�ʤ񾭖����y1���K�8;�Dkd�k�%+^�
��-�K����h�l��;��'�r�y�&��w��i�Q�vM��HA6�y	͝Z��}Zz'ٳ�����B�n	"U���Q�X,H��,�p�𡯺�����L>�đ��w���%k��'�3�k�%�`�kGEד��ib�5vL�i�mA�|�<�lEʇs��#�@��wr�7��4\�ﶷ��YkUB#M�}�j2�|��>�x�j��qْ&������:�o����^z�7�9�U�p��� 1Q��{�D1���W'��	��H����
y4���ЬB��Z�9�l����D�=�1����hƻ��Cɨl��/(�����I���kv5��=L���-��ϰ�R^Ἅ�Sk�L"�	���v0�X�3�J-!�A���|$���vj��I��V�l�L�Y�oג|<�'��>i�j/)�'��;�}#�#�SO�oF�	{h��*Z�l� 1�����S1,PT�|=�'<��8�D�Y�(嫏�'��da��0h�ntɦ�2�-
��)x ��b�o��>Pl���t��� ��HD���w�G[�0��SB�K��QB�C���m�;N��)�4���Ybk�H���!����储��
��rڼ�QV@[��!y\r��Z�׻�/4n��9����f���r��h���D�9��E�������tcQ�U����X�]�/������M�G�Ο~�fM��i��C�lY?��sX�*]��5�9|!��tb�Y["O�6����v�+jE��J��{i�"�n��_��1�#�"�[b#Ql���ɩ���ɢ�Q)��)}@ݦ�Ücf�Q��q�'�`e���o��w�t8b)��@�/;�r�	V����Jon�	*/�ק��S��~a|���G����xd�Iu��xt,��d�e��@o�{S��;<Q9V����u���.\��=�dg�(� ��b\.�������d���ڵfH��Պ�K�8�w��i��rڳ���sG4C太�f"�W�k��`7;���ٮ
Bփ~�����Q�"���| �D���M�|�=0�Q��1���\U�+�9�(kCɿ��
�v�T~
#���@\[����dz����d������B�T�4@����ñ٧v�r�j]٦�LeK
�R�n�[mXvEaOjj�m}
� �Ռ�6��/ԗr����	{?�19LF׷�qj���Z���_ﵟB�Kܙ��P.�l\�P&m)��҆����p���=�?����?�u���Ę ?��B�~�2u#�� ��r�k�^Ҙ���q�ѶP��u�׬c��4�=�M=�x@!he+���4�'�o*KvD�O]?���u{W���d̚8h��a &���GU�S_���de�h�wג{v�#�{��&���[��'{��&+�ˎ�.���V?<I��e� ����9����J��e��i��l'�!-xS'��Z��Wȃ��Xgi܏]�����W��u�qB�^���";({���^�8t�*m��������Ȍv
I�#z��Ș�0ʞ��m�ȶsU<,�o��H���|>�\�E΍d<�փI7ۉ�\�\�j�o��--����t[���vr�b�d��ԑ�RQ,�Y�- NS�OO���^��+�l\�',�wl����n�@^���>�3��<�wм�ܺ�2sm8��rek��[*�UQ�K?,p��e�F�arTz�Y�<i=;m����T�9�+e�u����Hd?مhBHYY���;pǬ
7G���go�@�n.$6��<��Q��s�Y<��ɚl�%��y*��A� �q���N�D�(<w���Yh��}d_���|`���igE�4M�/'�_Rn:��ވ� �;�����^��1S�"�v��*ߘ3;l9�l�[��u�#@�1�g�
F�K���ݿ�h�N�h�����_�I���O��.���e]��{JH�v�_�ĘY��Gi&;IzΆ!�j��?�����9ir18��E#�'��z�Ȅ
�.�#$W���?��g��8?`���R?�|�k�p���ڱ�Nl:�"W�w�J!�1Ϯ�e��J$X�9��
S��X��Ii]��!�����2Zu�
N1�k��%���r`�L�ʟ��&���&��=m9�,{��zq�R�e�1�~n�������#z)�DDL��Ã�-�����u�����Ma#��M��77@��ri����/PЀ^+�/��r��4�B�͉�b9Y�Wԧe��<X���J��CZ����E���fd��ͯV�1^m�P�&�C�n��jwt��Uo���I�#^	�Ŝ<y����`�*y����7��U���G�Z��D֚�$����y�
?9bS099��H�e=� 3i�.T]�����5�`�1�1�b���G!�hT��&��޶�h �u������t+{X-�v���#�aɫ�������k/�:-#5�J���H�M���L�}���[4;>���?z���E���^'���K�CJe��>���� T��HL���c���͂��'AJ�a~�rW����EBOnoq;t�����X"��U�z7��"���;���`=�)?�q]6��RP;�V&>N���@�&�JC����/�SN��ʓ��xMI|!�d�g�y�Y3m㲊��]�Sk��x<ˬ�r��@�G���fE5���L'�Y$�R�2~c�����^�8X�[_軋d'�'�);��$[�R��7iT�p�.�|>&Z,�C��(�K�CAnS�Wdֽ��!��LQ�c\���zT�ݢ�ė�@b����Zt`�n$Tss�1;�m�9�G��9�᠊��_/J4{��Q�fX��r_��0|��5x��W�G@��A�Hᱻ�Rl����h�]��\���Mr]���ғ*�"\ǩZ�.��ۭ#�A�)�2�`%u���+�������"=x�c�h����^/�qϑ&�<#Qt���"�O����=@�竦�+�=-rƨ4�h�s�9���$ͣ�W��_a��d�N�y;�:��I�O��S��H2db������a���%-�X����`�C"�9^��͟y�d�ֺ]��I)c�ql����/�. ����j�\^Q�$�:���L�o0�����ĈL�	�ϗRc5���|ލo�.
bV�?K��BL�q_@0+X��|y:�g6���٨J���Ж����B�%��9j� u>o�m9��
rA���>�	���+"3�A�����QFÙE6�M��sH�\#noa�Ga�K�m�U��W�m	��q�����3����Q@�$�԰��M.�j�Ƀ��ß�u��q���}�+lݹ$&7� h@o�,�?�~��Ki���\��&���nC��O�ǜ:�z1���S�� ���[�H��uL��PU
���������Tx��0��v-������#��ت�ϑQU~����2E�� G�J�����:?x1���\T�R���H�l_��آ\���F׉G�<�iV��~ou�0O�n!mP��K�8�F��Q��J6��>j�?����O�PP �!�������c�c�S��O�,%�r�[+��/x���R
���Z]��	��H�7�����W���y������a��qP��zI4����9'����W`@{9,�[
��J߳�m#�ǻ�w�M�_�h���w��;I�+:���P�h �zЌ����xgԨH�6n�"��#Ђ�nIxӔCs!#��r�����2���y�tK�0���H���u���L^O=fP^�ղ��|z,���+~�n���:�z��/�d��t�i&�J?�b:�KC΁��%�\p�)!e>$��O�(��R$gV�G%�tt�X���{O���qU^Q�I�OC�>#

H��c�m$�Y,(�UDq`k�n�\� ��ZW���"�a/<�u	�:B�5;$<է�~S�ȹMX�݆���_��h�l}'
�Zi�)�����X("�Eܤ/}Y�Ex5�Sp�~�%�%�xOk|a����K2���k�yfn��vq^ǥ'��ZN�<�l��Ru�If����s�G%"�������0&Jq>�N{�ɗ-�Rd[����"�#Ȟ�
�9��1�~[�0,�jN�m���9Y�� z�L� Xpmoplc�a@����c��'=;k8V=�F(&�!	��g�����|�V����W�y�jw�d�-�Y��.�Y�mss-?o=>Og�a�{4ڄI�K��"��4��3�(����o�\�kD��)�~����l0U2I2�p��_ӟ\KJ�D��H��d��׻=��ϓ�����l�$�򀚴?8�*�iu�*�*�iӰՌf �˖g�����|8���^^W/�0dj��2K�^�ݩc�tȅ���ۿ�^z�n��7jԴ�����v9�t�X[���'�V��i9�'Њ��{�w��Q�T�k868X�x�eE�ײx!��l0Am�G�l�ugo�Ǧ��}>����x��N�r��~��#|�Q�Q<�����v���Z�T��ΆFC�O�b�8>!��I3f� ��l��t�vgyd,�|��yޣ���Y]Е���Sp=~��,�ق�d�?��؏ ��<�c���b{N�Oʗ�5�0m��@��8��h���+6���꼰T���E�@�L��z��_�Xv����ļ��0���Y�X���C֘Wk+$osq�P��U��鈢��K�g��?o��C��c���SF#TюS�ܓ��}j���s���#Y��Y $�����OW8��g�̳�=����!��>�����[e^Q�Y�S�&7tpG{��"ү���	b~.��O�Ն�i�ЋL��gmM��,�b�l��c���_�fh�:m%�=P��͚��U�^uSzT$M,-��-��^,��p��a�Qޯ�q�$J� t�_�#�0�M�����ܪP�=���T�J�=R%_iB�>C��k>���<pī/�s7U=���!Q:z�&��V�;}��S�
.ь����Z�`�u�.�e�B�)jLf8}�	�Ȕ$e�|��[i���I��I �`���� ��-���N�pmu�>�uU�pU�g�B>*^,y9�"Ժk8 �o�J�nu�/�Ї�'+�;�F4u�k��L"��w�M��}-�M��Lg�F�cu�L�����yQ�_-ů�֣X�6lF�fҷs-��8|o�e��Q�e�\z������ح������7-/��( ��_z�Iձ��j;�@�ǡ����RWj�+]0��������k�<�km����sԂ�#���6�l��,��㯠�^�>~�i�L��g�c���ynC��x�����q��|�9�DUc}[#���X;T-l�*Y&mU�F�ܷ<�Ω˯m�6a��S^	.R{�ɦ�A��`�Ya�q�5ZW)F<T���l3G���'���Y���o	�ӉI��$���,4&x �������R��^��fU{�zq����u�%ՠrM��x�o�q�W�I.?�\k��R��V[��gt E���ۚ�<��&�c�S�)��R��/�Z��#� [5��jB4�*`���kS�\��W+r��L�7��m���W�>5��������l�i��/L�朐�DZf.th
�7�v��u�K�=n�l
�ŕ��3�LΖ�֪94`�1*���������O��E������IՓ19_A�9��UùJ�:��Pn1lj�R�,����IL����;s��X�h��'_2.���M�I�| P�U�2Gk��u -Z����dG8�/¸Y�i���#�DO��yZ�G7!�a Sq��bΦ}v��$Oi���VNAò�6�/��Sv�~�s����^�$e��G���M�d>��n���8>h��ƭ�z|Ό���#rNN�������<�d�Rmԗ��j+z� DA]j���D��Rkn�=�AA���@Q3^�c�8��s��r���cz�*�'[?r�(Ė�÷ѫ���4LZ�OyzN(�g%��l�:%i�o�3^|o���yޖ���¥�6���V^4*O�-}�B��iP�m�1�DC�^lF�s��[�����U���f��>�v{z����l� |��D��,e���#<���C�I�����7Ȝjɖ�ɪ��?~j�t|��T`t�)�q8�Y�#pk����� B��?���ҝ�5����k�s�8Ə�xzS�+Y��7gM���/��-�	�< �v���
ߥ9�|lZf��!��ו� N�H��r��6K�k����d��eז��A�I�p���c\ǏHJw�T��k������/�  ��s$R �hJɯl���ɳ3s e��``{���h/�=���װ�BW|1�@G�&͞^~���z����Y�j@t������C"4�%��W����-��X�2(���r�e���*��� G9���VLb�0I�*��md�l�uf�Zq���$B�5>�]�$.��!/�gv�?4�r&�E$D�D ښe	�u6ؙ�+�u�|C��M�|K`��@�^����ɡ1q�K�D-TY����?����"���f�/��`X�7;td����a���2l�����9wS�5�Q9Ì=�&�J��c*oX�\ǚh(�Z�����$[a�/YFN�W�T�^�u��XO���e5����n����WB�PSJ)����B��,�HI$H[���E�R�oiʲ�U�P�o�l�!	��B��'a\ah��� y�`�Y�#��'�WdbEW�gi�Ny��Li��I�>����"��J�6�j�_:*W*M|�&��)ڲ�̆S^�-!�%,H��u��R������&=?T`�57맿�ޔ! �TӦ^1���xaQ�c���u%���B�(���#r��C�a��׶j=�� ��3���&�����/��{��	<���n/�]�,X��)�?�v?��z�N�*A1���`SF�%��ʢ����B��i�����q�����.�5PQ8�,^q��=[�z�R&��e��,$��������CT5�-%��'�`�td��J���)�ew�̻;�A�rpτ�t6;��`�8��� �ys��f���gP��p�r� 6�~���һ�v���H1��6����n����4B؃`+��n�\����L�����T��×�[����-�#�rb��4��T�|riJI� n�̝L��aLgK���C��C�: 9o'0\�]���Sгұ��G���p���/Ȟ�4��X�),�FY�D�y��-}-���/�>Sp�:ccPrt�L�"��h4Q�C��鈓��m��I���eܤ�'��'�9�z�l�����>ԇ;�xEja����j��� C��� /é;�Ǔ�}��5f��2u��W6���Њ�F'{�9i9ҟ�:��+8�����"OYz�?΄m��0�(�S�P� Z��-x�7˪V�M<vD�n�(g+��E��h��en׆''3W��6�->L�ъI��i�Z�����*ɴ�a��a��������sc�2�����tC��B���R^��Qn�hP�e�~CTgd{9��_�g� �O��Z�l�p������G	W��n@�H�.��ҡ�jQ#KP����qk�mu�N)
��}�UGh��4Kܭ�6Y=_�#G�c�[���씾ɵ5-@p	��W�R_Ȑ>_�6�jy|�Q���IE^}n~!/G�C9�J-���}ğ�n<v"ӝX�#+� p�3P��P	��φ� y��U�Q�B����xH9��8�Ɔ[M�FN{'ׁ�By�j.v�\_�␀jCU�f%���h�Fu5}&V���-{�_�����n=�%�5+V�#		2���ΏZwV��-�/�W�˿<~��!�\}u�,|9���O���|���������eK�:?g�r<�QAA&�J6*S^D�H�G(��ķrB@~빙�d��e!��mH�g�fFRV!��8z�0�+����?pM��e<)J!#����tB���̳BZ��|�����O���8�u�p)J�,���'&��ʢ˞��u,�/:�W�f]���'7��8���c���j��{!L#�)O�
@Z@���{$��I�{,kT�����A}����k��v1:�L�Ls�X�0!F��MJfF�#�g��]�C2���U'[7��:�@���S��x�e�7��{]+� ���N�9�ێ�6m��!�ߺ96ǨF�5�%>�YA���K�+Y�������(U���=Z|M��'Jͽ�" �\�28�W�f\�jkXEh�#���Py�
�:�-[���6�*6n�$��Y���p�v��۴���\�%�~� G�\5`u��Rő��M&�������}oz�\�ZB���tV3�|Ր���Tz��?��ڨЈ�� n*%o����vL��P�58��ɷӇL$� ��[C�`�C��i4��֏�Ү=0��_��B���-�W]�D�ɽ�]��Ʃ�g�j��������l9Q��/i�#�RD��Q�偈���=���$
ݿ}K��Ƀ-"��Bcz��|�h�����ha���
��-�J-_^;8h�`��;d�(�})�lE�z�#69l��wk���ٺꁊ��1}���e������<�K��W��/ж�� ��a��s�:�ys�SB���� �QK�X�B]"s���9�>���#�E}����c�����b�7��Vk)q\��ƜP4�-S�aD�J��Zfо=x��Mt	@�v`*�������4d�>HO��}/@	j7�`̭�&��J�w�����:\�&�hť�ށ�~�Q�����2��i?0Y�Q/���}2���<7��1�3޶��l��Uù� ��>s_G�G��%� �,���Mk�h\b��í�0u��澾�?�1�G�^���9���ZZ�-$D>���1ɚ�Ю@1`)���o=*4�ь�����aȣ�3�*W׺ԿԈF.�ܸ�|f��f.���k�ě>Q~F�=���"P#�*եd���˸��iV��[B�M��x�&F�דCm�~��H���iv��cO������'���pK�G`C�ֺϝ��ğ
����	_	����I�P�"�w�9�t�';��Fn��c����J8��� ���>��<QF�4�!�9ݻ�5e槠��*pssB�wXkr��齯����D���+�x�̽%	i�ޕ39��>�N��\0ETF>�Ln��l-�ݔ`����FՉ.hN��v��pK�ʢ	{�bۊrU���T����� �� G�#:��j1�jQ�_�p�$yǉ�����\t-//���,&�-�u�`穆G�������+��$nҋ)0��w@��d��qp]4�k5pmA�<z&m�P�Z���u�����%�R�JSS�����;��oۿ<���|���3O���R�W���D�����t��SQ5�`��+�L���������� Z\�&�]Fbm��݃���j�?YŶ�.{+����.F�,���[��-��zPAM���ܨ�?v.�F@�i��N�wZ!�$?OxԎ�h���w��Y�WE�C�ם�	�������(Y6�	1}L
����v�8�C����Į��֫��B�d���į@�tR���D����s��dX���h�����v^GvY�%*���P��d��E�	e����1�H����QÊ�nV|ƉN��|����Ex�Ȃ�⨚�=�����*E(#��.�_�L�J�(NB1�U�������8@�D�2�ؓCv�Y�ԇ�}#�>b<;e�}������c��Y��6e�8eyO�1�*�h�d�3j�!�o!&/{��TX�5ě�2�������>ׇ��*ԥ=#���Fb�9�=;���B2<����O���k{��F�ɋh >�3k�d(���s��w���w�Io:��X��|��3�|�9���Ή�T��f�Ck���}.�8�ry�]��A�mU3����)}��t:ydvU��2��)1�a@��"�y��а!<m��6�g���0�M�<(�ȧ`�q6T��b��c=�n���ܷmϊ�=��#82v��n��	���/��Y;',�78T�&����`]JG�+s� ��H�ᣊ��#�\`�ř��`>��6��6LC8���l��7
�"qq/`��0���~P��,8�@tc�g]�T�bS����RM����t�Q��
�%K(���������H�b�x���ZD����'����9��g�v�=�ΣNM�i&_��eN蕧��t8+۪�,�P�w�;�<�E���$Q:tŤH�dkiH���ʈ�ɚA=E�w���.���d�����}��;�'ǎ4��P�ss]\WyۺHo1GJ��XQDF6_r~!fl��		)O~uR ff=(q,H�aE�y?�	�Bh֓Nm��j���"�5�$�Q.��9+C.�u��໬�����~F mo����X�&_3XD^ԥ�$�e��7�闙M
E2|�1ܪk�v�1���s�K:'4��}T},E�x� �_,/��[�{�d�q�����6+ ���CC��AVtMYF�l� �Js{̚�ek$��8���Ox�~���]=H77�sk:m��ns x�-�1+�����^fg��x�S0�sD��9�ؤ��N{_�9%�uc���8B
��������i}�8P&WИ;�__�#�w��k*���:ضz-���g)�u�-/��O��f]��b���^�@�����b�Q�K���<1٣��0�J�:̧�Ѽ �,�nN?+pʧ� �64R\
�)á���5XumQ)�'��@��뀂�Aks��pv���UO ���:X#q�	��ߒC� X7]<d�5��T��Ӟ' �͋Ǉ����:�!D��B�w��V<�dN���QXłQ ��.n���F�Gp�Y��}�Oىb�۝�ۿņFA9\ش%��AҢ��&K��eyI<�aa�gU��" E� �ZBݼ=���������'�`p�fk՝զ@��Tb����:t+�lD~�=��)..��R�"
9�V��GD̪�,������g���ٹO-�`�|��n3;�Š��yZ8����-h��KJ�߼�����!��;*;�ha��I��"�n�Ж�����5�B�sU�&YԒR�joQ��/)GGȍlj��0�BY�QU%Bś�p��&�כ&�;�d����V���ca�|fFG9;���0��Y�Â�x؝�d@�Et�����%p�DWh�׽�Gq���9��r冊j�AFe<�������F�$��N���{iZJ`�LS˜�s�w3��;��A���u48o�h_���P�,κ�vN�&��eid�;���i��"m-9�Q�j�:��-�/X��L�G`�5�G�%�M+D�aJ��f��D��|;5 L͈���5gɏ�8Ч���	Z`�����V�K�d�u_�W:Rܫ�=d�侹��]R��n	�5uQ��Yϊ̈́�V#R�vKbtzna&��l�zM������)W��Q�%�[	ݚ��4&X����22�~ўЯ��G�n�Oh/��&��*M��y��)T4���?4jF�]
B|�i���T�O9���r,�3�Mn�9,a"#����j1=�i��(:t쏣S$2����!�
}7�S3��blLa�B� �]��jT'z�V��5_�?K(�kVv�뜞_����BQ��p��%؀\��憵��v�i�F�����\��>�����<��^��Gh�g��Ò%�Tz0����.�	u�����V܃�� KYCD�]�_�<��Jr3��Tx��s��.��ݘ^�<�l�5ݻ��s�++����`=�{6�w0CK�y����.�z����F�Ŏ�Q�s���^�;�D7ݎ���9� VW���њ�S���7��j	��F�k�	�e��f�_r��~�2�ᓻ��\��.f�O��4Q���Yg����M��żh^9��������!���]7m<��I.�u@
k�$��7�\������.����� ��e5�l��Wr�������$�O4b��,x��oB�&@��ȭ�y���m���8�Ο�T�>�8�U�s�;čo����
�̘��޾��bx��'/u�����4��[zK|���pt�K���4r�Lgڝ�UǨaiyK��q�0/}7���:K��.T9�K�+���9�@�����k��gQK�9�:R��b[b�D�%�z�K�@oL*�X-�k؉˙c�^U-�gt֒�~�694
Ѧ�B�):�i�v��H��jj�S�xX%gP�c��j�-����[^�3��� ?H���	�.S=.jҔ��$a%g���@� 
s�T'z�#ۚ�u3�s�o�=��%���!��:��Yԋ�4���˶ς)^��2ҭq{ݠ��a,9}ЙA ��p ��Z]�;�����<.au�1c�=[�d�{*�q�GV��Ek`�ٗ��?<Z����Ak�{����u�-L��'%4]��E4�$vW���e�Yiڛ�5�#����+�.�HRx�A�^��,�N�Z����+Nέ?����&�LX�r<ś��F�f�h]����)�ܪhr$�a(
���4,�+Bcϓ�Bݧ`Q4��X�Z�𓌅�y/M�M��<Gn5�0Pd}�DA�BE����������E�ʺu�!�;�E�O6�b����n������Z���y��q_u���P	�(�M��9c����xϤ�.�9�dþ%"N�J��1	�9A轒���O���b��@���%ER�dj�Nڗ��#�9d�bbSg��g��Q_w��������ˀV:���;�GL%R�Y�5m_"������}��Ȉ���tp�x��I3���C���o�E4W��;=LsP?5U���~-��m��ퟘ��`7��!(��W����}(o���i��q���eGmϓ�s�@�A;k�C"G.o����s���>߾���&ԛ����*YR�3̰]��6fc�N/�����%��&'w|`j�
򿋪�K��}Q�S����R�t��jsHGK�M�_��̢��	�+�vZ��#<�݀\lD��+�p�7��inba(�nW-���f���x��'��FM��D(I6
&y���*���6K�U(��O�w�Lɜ��z�<Ed�qO;�4�a��9���_��2���)���"	o_}S]���-��m'�b�T�&���0_~(})+�(���B�g'�?��1�4���T��Z	d�'DB�
K;��6{���C���:���!�&(�5��a���H�m]���MC����#qԵ�j,�4_��[�ܙ:v�Mɮ�䳳5�e��n��%��O�M)��vo��6M��g�����,`���������-"���ؘ�6�qs.Ds��b���d�i�J�",�%��<�(�J�b��Dm�G�X�=y����}qJ��m�&jLRW�7'�&,t��Ǝ��{.kS�qI^{�ty�f��2 ��.¨�s����<o���Jn\�
�<~<����Z�$���/|�[�� �5>��1�^���@��)��]�v�dC�Λ�4�`�����{-EP<�<�"�������6>2x�P=z�ZK�Ąjk�b��5��� JLW��ka����'�FZ�-�}��Z����F�Rr/b��3�3���t�Y������g�R!Y�1R��4�_�(����n0�u]X��ڑ4��&�W*�4'E�{�F�L���])v�iAܭ�Y�0�t����L�/@��RK��uL-��#�n�rN�Iq"D	?|�s�jU�q���NV�>�"� �i����Y���EdI��2*��L��/�eq��>�j-쵼�ܡ�i�a��7�f	�N�P�3�2�_COF�:�f���K҂�%�)F��UM��Y�^�d�e������@>$O4��Qw�.>�پ	����L1����n�h�V��4	TyA����i����/�F"^�Ǔx�4&/��|U˴5{��	(
�Z�3��o��|^Fu �.��e��D"X�qy����9������` 4n�}d��)���z�J������U:ڊ�/,��9������7�Q�0VK�ԴsN`o�T�pW��p#�5%��x���������o��E����0oFpB���^l�u�eʀeR݀ʅ�bziZ�%b����u|w] ]��+
�_/�7������&~Ӽ`���X܎J
U2D����ֻ�C?=Q�,�0��S�bO���=z>�EB�a�x(�0;����{��y'#'��}�14�V5�����y��:d�b6���gÙ��U>ś�E1���i'�p8^��$�����@%�T�6 ~��_����%�P�޺�v�w�]�;Y�P��`@8�?�WBhVEG�u�z��,�۾���:_�(H�~����l�Dix3��x`���rA�3�i�������N��<k ?@.	���1<�U��^jK�u&��6%��Y3�R�8y�g#��6��E��N����h���(~�A/���Ne�ّ�:�̂Neߨ7���1���15[O�'�V��i8�*k����:n�F*e��$�2�#��ɜ��8p�T�.��E?���J1_�N��5��fo~3����8|�6eBn��/J�H� |���Y(���}��x@�#�S],<[���)��	�"�&H�k�a�)/_�p8d�͏�L7O�Lȷ����G�U�?;
׋���3��W���q�Jb.'�9��wL�J& �����R���}y�ys�ߛ]�KaNv����:9���n�7�3ST ӇP��h��r�ʌ+V'2����S��teLyL�m�`��Vo�qE������˺[v��p�4�n�tǘ�Y(mVd�O���E�M�]�{5��Ķl�k#��0
	��'�O�R6��|����f֗��Z�r��w��Ũ���T�a#=�D���\��3��J�D��r�Ǫ���l=��u6�"�&�`�X�k�۔P5��Ο�{�?Ē�Gu�;n���o��CC~l�y�5���<�P�c�S�ٕ`묩U�1��\ʆ�;�BK7yd	C6ޢE�	��QM*+����6�~�k�8O\v^�9O9�؛rp��9���#> s 洺�P�����g���7Uр�yA��R�]ȓ>xޫXA�tיb?�9F���0��R9 ����ۚ�]?��������0�*�R3�m��{Tr��+ C�~TL��༹��r��ڑ�VI�F�8���ͤ�X,m �Dr���,	&p�����������C�)'RI��K��8��<B����SVۆ�����I��0zl�]���9��#E����'���4���M�M�\bI]��T̜��$�h��z>�����m�i�k�	�i�3N��%�4T=��dyȌ��y]�B㤫<�g�W2��^	�B�����<)�g��:�iTi�~�6c6��]���~���;���k�5�]�ʂ�e �
�j�1h��n���q���u��l�Y����PZ4"p���f(�E�y"�,��3�k�eK��.�� �	y���xT6�J�Cs2>}FB���HY/-gƁ��7�T���n+�J������;���ycE�E� /�d?�r<���4#��r ��^���GyAk6����e���.� 
�ԛ%I���I>�&"?��D��n��l7ɖE���ؽ��	\�*ژ&O`QE�2��]a�"��R�c�2��2�c�V\D��$��]
�M�W����2�l�3`�}̱t)��		M���`h��KU[���G@�Ĥϟr�9�0.�LdƊ��f���7rQ-�TZ��4�r[�F�����Oמ��1��,�:v�kև�A� r�����O<��+T�C��뛥�z�����G�f ];/�;��Y#ϰR䓩�"�-E���f�����o?�{!�uĘf�xFVq xf����5݇ǃ��s���k�T�&My=��_n5�����'rA�4[��F��@�gc�ǌ,�1�h�����&�\�F�c<2��`D_�r��(Ŋs��#�HO�F���!l�g+��й/v��S�к�҉��f:�2v��R��=�������%����v7!)ጬ��1�f��Sly�f��(�t�Zsʣ��2#A I}یB뀶UF���'i���d���G[B	�dAւC�-�ӏ~0h�yh)�e�R��GL�5dQ
&)���tuT�*8�9s��c���4���Z��.����[� �]��.��!�9i'@���-r�]�_�u�<�E0�0�����3w�ɴ������>��*�9|S-z�����6P'f����W�J3r�,�������w��dW6�B��X�@_Zh�|�Ɛ�Y=Dţ���%Z��p�]P:eVmz�U�)?�ߔu�S>�˧E�1��v�$�XJ	�	�V�|N�����6g�2���/�6Q��W@�� F�(X��#/�A�O(�TsE�+����G�<;ޙϹS�Xbܘ3X�!��祳�Uf��2pxf�\>l�Uw<c��NGdc�����GI%E����[����.X@�!��:��Px(zU��gF7hu���+��r�B0�jw�7*���.�]�{�Α�A�d �g8�XUذDj�BH�x;�k�#��4;�Yg�W�c�a�X/i	��Oxv�ak�B�j5 �z8�w���S���  t$����m��N��Q��<s)�D��	B�W�<F}Z!�lJ���l���H���bj�:�oGN�H�[��q��U�O�C	�l��'�����u�<�`J3�@J�^�q��$�I���^��EU� 8�P�g�l�T�dhY���g#��v=�_������7g}&���G�E3F]���^�gܾ/	J��F�'n��E,�R��8^T��h6鰐w�ժ�D�*F�6Q�Y��ګ�43L"!�B<�E�߹񿆜��V���K�}�2܏b�[���u���iw�u,�[t��R������ o���@^�j7뷟Dq������?��m<�nr1�
z�}Y�^�t漳M�X�aeŨ�gK��.�P�6\��T�>jlL{�[��rB���1�K�o	I�d�5п�(`�|1X�h�@R����>s=�2\�:,��^��ǂ�:�Y��|(��3!K#͌|�OJ���VO�r���n�9:�W� 8�k��{=�s�ͼ���;<	-�OZy�6�x��e�?�(A+|���8G�Q̫�9�E�͔��<��jZ"P�"֒-����B�u��lI�����Q�����E�"�q[�=�7��V��x[K���'�es`��u�K� �&��c<��C�ItO��U�ˡd�φ�M���yk�����߅��{-���;�)��I{z��R>fM�}���C
�8�_��Pl��,���D�1YwsTʃ�\?��m擽����D�N�5������Z/�^��BEw��iл���-�&�o��M�.� �v�q�/��h_�-��n� S���<�Z��~^�3!!���C���
�������߮��3>�5���|�����|�;���}�j	~V�ǫq�@/aƽ�����\+h%-��[��W�vX���32�Z�p����D�:А78�x�@#ׄe8�7�bt�/}�YQ1g�ڀ��L׏[���z�1L�Gvf�D�?� J7��K<Y��=0���VU�{�]:�o������u�{D*S^�a�u׮q�͑��vC��F1*���]%\�p��: 1�qIĭ�Z� ���k� c38}��;�\��T�ξ{`F�u����Y0y��<a���񅗍�ƹ8�2}�)Y?)r��D��8��݊��SAD��yޓ�M�>Ps����A���vt94�1�� �gK�q����Vb�9UX�U���q���0 �A.0{�R�Z��� ~�_q�zk����"AA�Q�S��� �Y�77T���w��V������&SW��o�`|���`�|q���Ǔ`�#^��z]\I�� ��S��r�W�-jK_ɓ�����9E���V��]"���e!g;c�)c&�����nk,��ý��$!�-G�9��#m��ĥ��u_��z�y��s��D���7#�?��pk��^���;}��u��+�F��ϳYRf�V�x����E��u.��״N�H�.�R�ՀP U��|�P�13�A���N�UlF�(R�O��Zy3A���WL� /'�L�3�5�,�hq�hI�B����7�$��1�X�MK�4_񸐖~5��%��������hC�X�b���B7���y����Yf���'�,�� 5P�δD{�G0�����$�$��5.l����*��,��IǍK��*՞=W�� a?!��S!-���oV��(v ^�d)�,���fj�<_��s�:Ϙ+�0tE����8�/aصBx���ӧ�dk�@Hy&d�B
ɎCsV�ӄ>���of������ɘ�f�d������{Mg�[A�0�_F�����f	���>}Ui�����e&f`����h���+��r,�ݮiw�cd�h�?���R<�b��PRI�ԥ�N�r��mD�x���2M3(������m؏6#�\�~�c�k����)ѡs�x){_�İ�E˖��W�ڦ3 �Dhw����c.�N�-%9o�`I�V���N�rII���`�(O��8��B����P�YBE�!'8A-�[�lU�J�Sp�ZKB�u��٧�2+��D#��U�=z��AI��)���C��(�F����)|j�r������wjצ
Şx����_�:)&<0�'���E�`+�V��@o�ݫ�R���4�wp����[�lA
�B�Za�$ZC�
��YFq����Ӛm��\���{m�9J�7���a���0J,]L3�b�&��q�RKȋ���vEޗQyj�c�-��$�n8�?�$�JO@}i��-{m���`���%b����c�L>uv^ҐZ<=8�'0��.�����r��w�.�r�$4<?��!98�o�1G�.�&S^>���&��*̅ղl���`WO|�
��bE�h�~�+5��>A!u���0DB�A]Ey���+�P�9�\���_ͧ[e��`��|�/~`�Edr��~��n�ˀ��2�C8�;��$�Q
G%	Lq�F-������Q�9�f��'fTl���0<,~^~��j���"G��U��g�
%�l�.{gd�t(���v+sV���r�y�`ϖ�s}�
�W4��?�̊�X�ka?�l� �(Z���X��嵫�&�|��0����1�x�{�\X�-%	�07(�{�BĻ������b�2�b&a;0�!x�V,=@��Ƿ�$G�A��,4��\m���'Q25�9��.��7���ю?ӫ9&4��-�b�e&�=�����X�n����ɾ|��W$��#{)����b�zn����9�Kknd��'�Y�1Tu����H%���[��`5F����$�gW���3�=ZZ8�a��!�)Yz��)����͚��DX��J�l�Q�>n�W��CL�&�c���(�0�����=!��iOa����J4��]�&<.�O:�
9��D��s�����Q�1t�w�I��E��
�PB��U�+K��!е���c����񻄬=֮X�^�=|���~7|�ǝ>�q���_�%1�?;|80չ���En�DG��t̛\DO��⴪owR� ���Q�� �'"�^�$Cߓ9���/�u��=I~��g��p�[��"T����ҏ���z�H���j˰�����+oT�u ��@y�:�Q�_R���ز�����c��%�v���Bw��h�E��ʚ�rʲ ؂�:��3�.	sb�'B0�y�ef"	��+��?��}�[e��d0�x��^�$�S�a�����}��4���/���"3�uv �P痫�[�ѱL^�)bq5�����r�Ͱ��xE]1��4`��d�o�0Jya\Y�,PH��w���0��Rq���{��l���3A�.�s*�9�z���G�iW��;��Y$�q��A.ukZ1,?�a�z��8�@�ᙲH����