��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k����W�z�N��VXi^�p���d�����3X��#��*�4����^�B��os�;poX�Mv�Ľ�g���ܿ��q��o~9�c@c�s��i����xw����`""�G)W݁ꍘ��zaheC�.�)������f��iE�\x��j��X���9�ƹ*UW�Ƨ�[7H�I�����1Ԥk�c�+�_�Hú{kdm(��U���&�kw,��a]oD(�#����F��ѳ�m�-�F�G�ߨ���:�v@�g��=�[���\�<��.�;F��W��Kv�Q�?�;�w��W�U%Y5)_�',D�#~;� ��W�i�تeO����fx	q@
�+���`��Z`���4��j�v���`<͊�kO�Ц�@ȯ6��Ag��٧�;}ߑ�EK���`�:!�G�F�Cx�t�0���U��/�T��mmEC_O3�ј1�h���KCɣ^������DL���i��� �'�$q��d�T|�������jC׵�k2������*�3��4���h�Ґ�&��?�L��o�,�)�(�=�c���`+n?���*r"Y��lp��_�zA9#|���ot
seU�������i��@�=!Fֶ��mJ##���&x?��D��8�^Z�[����Pn�UY����#�ɶ�zi�+�
��
�m8����C�Q>�M��%�JS��p���	C�N_�G�Ի�c�/ʠk��ڥ upN������1��^O�3>Y)�f�6��dz�7��F�d>�h��^�y�%���.d��l���=�$R���AZ����o���4�e���|0�Ǆw�l���6_��3倪l�S���Χ�}kdx���)Sv��	��A�j�jM$�Q���v� �μ�MZ���JX|����(|oYٰK�Թ�*,l^�����dh)|��R��S7��_[�gU^�o�w�,�H�r�5P?.N��Z��c����,Mãl��Y��� y_��>��8{�����0�6:��%6k\!� ���iZ�k�د	��p͇
T6��8�&�c��X�I� x��F�f�^�4�h���~*��.�@������$�V�[/�_~�չHEX�[˸�7�J�]F�8��ϡ��∭���>��"�O��ō��F�7���k�9%v��Ge���$�Ѝ�JK]���QP;�S�@r�����*�\g��Bn�B�$������E�g��:$���/9�)H�^ ��i!6���ސho��z^�`��I�K����1�eh �D��A��"���,��[���80i�B7�E.���4;I"�s�{Ge��:��P��Y�T�o�B���Ȩ�f��s54��C�``�����]���-g��ܺ�v��q[ù���5�כ�-���P�O� � �Xb1e���:t*#[*B���㕶���b?t��
�� ލ��\O}ޮx�U�S�`X���v�Imu#�\=���4�>�������c)Y�9o��F��<�G�$�k�2�7�����^W��V��N"{����b]�
"r٘��?��D[x�z�*h�S��O�mz��U@D����zW��.4	_�ts�v��]���KoC��"ì߉��L��d�|�����e]Zy�s�B�5�)���zQ���Ł&+���Ff&^o�������U_�����٢ك�� 
g%�9i wT���)��,�֭���t���*�.%�5'Ԙ�'U5��i br�z�cOWEZ�RC�^���$C/�z��;m��@	INq'4��*+�اtɼ�N�[N6��"�!k����z�%93Z��Y���¸�ӹ����q?��&p�Qa-q�v��fn7����V�q���N�C�������N.Abq��4R�R��86ᓣ�w�p�+���v��ʢ7�KI�aI2�,�B�?+����nsřW^���n�\E����{��.�ygfHZ̹�F������lJ�u��A��������5��b�̡I�<��&�4J�����z��@�e��������4�x|)��X��q�e~��鑶R��+J%M���{E��p+,P=��͛�vg�KN�g��b��z��ORh-��_^k>#���i�-P%d�B)��8�AU;'�*`N�mʿ���kyL�aM�k� ��Pbl��ٌl�7�����i�)zko�?�N����ܥF�g�t��Ã��5�=o�
_����!(,8�M�u�7|�PE[ƈ"�X�L�7�?B)��ֆx��� �w��hE4�����D�"��+��h��B;�m�٢�
-�����z?	���%����e���p�*����̬��z�|@��l��
���p��V�>�u�h|��d�NJ�=8�v�	h��㝑��X\���fx���π<�	}��P����������q%򥉵mB">`y�'H0�k���̕=�� ����|���BA>�)���D�pб��&�gsɾ�Vʘ�f�U���nJ$8Xq���d����;ͺ�8�W�Ĺ���J�XT>��ۑ`8-��λ-�P��/��W�UFx7>#�b����G���Pi�_����*�8�����+���ʷy�m/�D7YuI�H������[�� >ٔ* 9.2Q\��3=���##Y���!��ě�����;UrU�>�{�����$m7�pJ����������E�=�P�f+�3�3+U
0q��'n��V?��� â�cP�	�o���elI��b�:���EƆ:�VA��~O�1��[y��6�	?�[�o�!jHe��\�ҹ՘d��=��}qp�&�hZ���g���A�M���Irl��3���~�T��0y���R����򙶇�9}e��chP{�{��1Ȅ�5D��%I{;x�dԥ�5��nA��h�,�Ip{���7WM��G&@�J�hR-Af�f��ڂ���h�i|ץ)���d�=�ZX�8��_"l�Ƙ�jɢ����<RO�?!��z �o� � ���%��;�raIiyja�EЛ�1���}��%��7�,(2�ꇷ�U��ߜ7���1��`̐N�B����b�?�cŖ�mmS��6@� e�oT�K���Aoi�޸�,�?f��}B���@��-d��Q�r�l����}� k��P�$ũ�]e��;����ʈ���T����)����S����f���G`�-j�z���@��1I�������V|0���Zu5�?ڃ0�7�@Y��r_J}��pH�^�-V����H�%#�������@�W�M�Mo���ޭ1JP�T�����ҫ�c�T�ZTsq��J�+�\��q&|X=���Yފ,_��x6ν���r��E>E)`Q��ɹAR >'n�q)(�;kwN(�>9�}���>���(�����)��p���7��MwR�C�f1��O>Ve������?�l]Jp����`+LE.�y�X�|W�P�s�5]w�'�:&N�;/�^�v�^�S�20��])&��Z;�� ���_��/���P�<���v~?�l?,=42�W6����Q4V���)���j�E�D��-s���*�7�g=T>V��y�w��p�	և�}����X����1�.}eTJG��C�W�詆sus��^�KG�s����b������,.��6x�S��	���2qFϙ�E�(���ݶ���MS��3N�>�A�Ֆ���y)l�=��^���	�}�f>𝃀(�Ɏ��U�nHW����1sH	~Fu���HJmf��Ov�*x,7ќc��<a�-hCa{�&�����5-v�<�ߍ����*���#z�m�w	j�����4F0��tx��DR��b!��W�����_�������D�,5��(~[�_�}��X��8�og����\�c�9�K�B��8'�{W%4��f[~|J ��ڳï�!oeDI��ChT�����K�
�����-�If'#e@T*z`�Z)֋*
Ef0�Zj�Mp�7��"h�ڑ���o��V�S,�2�'�_w�p�&J}�m�1�;1�c�&�?k݉����i�5`���P�3���V�'fd^E\���6��,�b�/��Z�̀��Gq�	:W�Ma/�57��sd6����YP���N϶)Hz�|�o	̙D����q��w"�d_<��E�FP�V�ϿHWړQ�9����)���[���}��D ��9�4��Ïw������jr���'qgL�-��ٹ'V7�C�Hl;.�����0b-"k*(c�4%��4��tb�w�25EE�/���0�oz&"kv�,�3K��ڤH۱j/�,���%|q�'�4�P��L���[6>^�
S���=���'�8��P��Ɔ��^Ҧ��H'KY�3Q3���!r�H�v�����j�V��^��E��$[�xv�!W�F97�Ur�����n�~:�w�AQ�Ƒ�b���2��qm�_���55�\�hc[*sM�����{-���8���4���k��y>�Xf+��%Ɨ��ˋ���@��W�9�l��r-�݋�ִU�m3�#^Y.4�����g�񦬡 	���R T 4�R��]�.�x�,���C�#���o�b/fPI����"��)zҖ|M\}0�s��O�B8
"D>�Kz,��P�s7�^5!J��0��⍼-�~ ��[�_9�jÊ"G� k����D�o�n|T{]�PojO̢8��ɏQZ+.>�>@�N�n�e�s��M����ŷ<R����Ϭ��kd@�=s�@��\�=�cb��g�~f�䬃t.4��$��1���m p��|��^��j ;d�7w�f��@����ͮ�4C�؂��WԊV;��K��Da�Tiq˳H�E�lW(�HH��o�6�]c�4A�&�oiyJ��$�f���(`1��֞��2vc�ZE���	9�D�q��2�zu���_��=��e:�?Y�Ћ���O���TN�ɖ$v�y]�@�F�T\� ��kX�c�6k������6$c�G�씶=��P�`}P5Q��(ɚ&ҽ5L�^��gF�Qu�� ���Y�<�T����L!�{�iH4Afa��3Ť�>�Q%#����P���=&I� ��ff�E���W��YR�v��:�6c+�,�olJ�I��O��?Z�?��9�l��o�����Ly,ο"�}�	{I�\DZ���Rp*V�����ǫS[s��Z�����{�kqU�����	j�0	~�ime�:@9�,˕�C�!U)5��>sh�����>�?6��-|��`!z^���^��c��%�q��ǽ6�<<G��O�9�m�r�����G�`����8Gv=�L��eL}�J^a�lh���0�L�2=��u��P����w4�jޭs.�T�_KEˍ����7nP6��Ws�=O�E��~���jaf=]����� �c9�@h����n*�;>fӶ���!�A���m���U
���?�7K�� H]��3�v��;�$�	.n�7�ɟT "���0w�lȕf�D���G(�L{��iN�L.��,~�d�fZ0�FQ��IǾ�Ba�����d�v������uJ�- ��%z�F+�m.��?�snK�DB��ڂҢc?[LsAL��D
yIxՃ�=�% c�]��a ��
-�z�x�����=Ht����ޯcP��*�OR�hD�:�n���~1�r�0��׭��7=�����&ٖ���QʟP�\����331;p񔛙��
�K�P��[��*��	W<�� !}8"kZ�ڠu������8�H!��S/�t%�&.��U�Ղ�9�������CX�q����:�D��;Κ(*g�Jl̴��TX��[�����S�?X:�g�+g������"_�"]M�!����񦈳�6<vR��{��	c�����a~��������d=Q�ؤ�+����լO���FEz���d6$����ť��5�ӑx{V����lk٪)|�e�L�1AMe<��#]Vdc[�,�6x����b-���
��v0�ꏁ����_�Me�3���m�=��KUf�7�06=}�t��t�y{�|�� ���*�Ud2�Z�=s5_�6�2�Z�m��0r0?��ˢ�
d�W�PT�w�O��e!��n����i�uW�����M��ʍ�����:B�h5�z�s�(�K�4��g���nI	�Ԕ��囯�xNć�0�U<�I/��x�v!�,�<ﻗ�=����L�z��6.�d&�?j��<�*��L�Wx\��ֆ� �Ta|:�v3ҹ4!�:�6>��F�环�����B�� A�Ğ{���6+pė��b�t�L�'����)
3�$�SU��<�Y��xem�Y����^���\&����x��ej�	��z'i(#�~s'wC۪�Q ��Q����f�fLp�F��g��2�:	}�=�M	�M9Q�ϫox7��;�G9�~�Ad��BF7��<<���ڣ��kPP�LR��
B��1y;�&قJ}�ze����d�"(@P���8�/TB? �y�s$q������P���k�V<(ˡ�I���9��Юa��Cg�Ӓ��BKڅ�D�(M^V;ڭd�w�W�U6Tk@z0�QM!�)��P�i�>D�o�g�W�q���!I8����5�����)^����!�$�s�c�Q�>̈́�g��ս3ǘ�Ȭ�ULa�. 6��v��6�.�v�8 ��L)_)�E�V��<=��D�?�2���	I�5�>�^�����W#V�K���u���/� fc����iQw�sd��E���0|�B�����{�����r(�-HΞ�X��Q��
MJ�N�c짻�>�5�db�����ĝ������b�X��C��o!��u�G�&�I�so�h|�����
q�� 2�* �O���Ac��z��Psn
9 ��]|�R������Ҝ[G����O����'0.�T��m�Ѯ�̞���P*	���P�[\�f�����yv{c�dg�KO�m���K7Q̹�Y�'T�
|^+�3��,��G��qE�
J8������8�ءE�`��#�׋$��5<���d�,Q�T�]�C_~�ˀ'L�[������([j���m�@�����5�q�,��}�3.�g�_��7y�����'���l�ZS��������m��ָ`��ovPoo%����4X�� ��	y઼�&�8��������1���ݒ� �X���pp�8/lB3JXBj��I�ݗ���f����Xu�̩��j=L����A���'Y���Q,O#2����t;.|pY|�n�ae���d���Pi5�M�����p{>L�6��}�JX�M��u��zh��6A:@m�k�@E�[M��ʄ<jx~��h�,c^3�D��)� (����iބ�-�5$��?��Yf�H�� �8������J3�=��@%.���g	Q�c"��c�i��Qm
��!����鞞#V�T�Ͽ��K��Cճ�W�'�����rjL���| Q�q2Ś�u=-H�����������«U5�1��nj��s`rF�d#0,!�}Bc]�8[�$!��i����bIu�@�x|�F�棕|R0'X��M�ƣ%�򜨾�aw �r�u�b7i�͎U}�~�;����!V\�ߋ�����ۇ6��X���Lbv�V�ޠ��@��ɓ�������H,� �H�|�sH����]T������V�a�>[ƞ[�G7��&߸Ԓ���J"B�9�P���C#�h��x����Y0��	�%]i�,���C\ |tԲ�(��bo�o�,��K(7�.˖��ԩ�7�E���c�=B�JY�A��wr�ʝB��w�w�^Bn����5^�u��Q[L{��K�:I�FV�4��62׳�~�k�vm�p�*�yA'�g)��}Ex�8�{
�^�J�'+w奔�7����{�$Bǋ�ƿ�.���n����@4����&�����U}0�B_�RƯ�#�C���4�ZA�:��Kh+ɴ�o��@ă�n����~G̓�튊Rr�2.͑Ē��noA�qp��~�~G�)$�q�t� e';x���3'+>�����!}�ULp�Nm�L"�ӹ�n�~����ʼZ��=}�z$������9X��U��9C�,<l�I��g_����q���<y��t���O@\167�v�<eM`^�c˭�\�1U��MZ��3�C�uv��s�8|̚�Jp<+� =���0��cPQ�}�w��Zӄk5�f7.���!��بl5&/���q� s_�h�%H\^&�{t��&�SBH�N1�#u��Zۉ�@�/��d;TF�{
FP��i��ZYP6q����(�p��*���ؗ�)O�	��(��B����<�g�OA�K�+�]�$��EG�0��@�K.T�A$\���ɻ��/ocS��OF`�V���e���D5�m�B3f��3�s;�\$%݅��S�8h��v� �D��!�gT,���6�"��su[�s���m(��u���g���/��+x����Z��E��7�e�c�N�7�o�5�S��y�v�c��ѕȫ[�Ԩ@� �!��U�F !�
���0���x�g%����\���uG18y�߭��R���~���ץmP��|ۢ����|M��;�h+2|�X�ɱ���|?���P����G�˄��&b�3��»�Q��>�v͵����*�r�M��;����	C�|�xi�[�|M�����-���H����0M�=�%����4�>�,��-裧7S��i�>�\�Mt�~���A X2�MO1\dy�S|� �O�x�� &#<�U\�:=qv�RǦi�邠gg��2ntKG5�Ĳ��*�oґ�$< ��~R�&g8g	[�܍/��a����榕6}b�2������֥�UT��	fHD�`}JݺH��%z�_N� � ��e��'�zK��@�"�RY������D���7#gWC������E�9�V�����-l��	Fہ�I��6�?vn0��UozbQH�����ѧ-�޸�Aja/f�v�9�ɇK����ҡ������:#"Q))cซ��aRa�3
=V�c<TP�ӫ�/-�@>�i��W"���*��ů
�n<��FAQ�ͫ���D$ۂq8�,�����4�����Ĳ���,��1L�������s1a{�,!Ʃ�C�棴Y�B9(q��?0𲱲Q;`e�./�([��kT�c����Vb�`�26����z%E e
�?�{$�l�j��ɾ]��y����}~M%��߆'�5oԴ
�9�/�-�sl4�p�O��Gw�1pӨ�s����'��@��S&!@�C	}��2.����M�a���Hq1���C�Ѡ�aGP��A���	�)UcR�"ֽ�i�]���vL�s2��i@�����:�k��A�l�"��[���]���t9>M�TO���þ�}��Y�Č��>��^|M��r�d��2��(�����t���1|ǩ�?�ޯ91�=�3����WMV����L4fglv��	,Ɂ���M�Ƨ���MM�@2�AK��������z���:���皝�\�7c�X[�o��<��	nA�n���3�鐫Ċ#$�m;��ͱ��V�Y�B@b���'}������U�<	i��Qw�	k�pQ�j�"�
����8ߵ�r.������S]�v�fg�'tFB�W���~I@Tr��?B�J�Ǔt�i���R0.�2c��I2H�<X�˺Hr�|��w�Z��#�f��?�p��Ʀs��	F��f/".��� �W���S�g�{n��[�@ͪ�fV���a)�ǚ��v�J�8H���˖���C�4��8	�/�	V|W[U����+��d��S��i�Rj�E�.҅�	�Ma��/�L�MXآ&Pl�W��-������3��l��j�B���
<`B�-�#�w�'y�˜�~�R�_�ס+p҃��ig��^�P�D�;!�A\~�����waf+i��L�����c����c��2F�l�3��`�Pm����ӗb7�8������Z:�����A����ŸF�M��pux(�ӭݦ�f���I'p�y�3����[j�@�¥W�3v�>/�W%�������RBn�%뱿��9�l��4^���>�&s�����2|. �p�F;zD�Ԗ��\�?��)��#����>�Z�����&�Ǣ�+9(��"|g璐	v<?�)&��:��j�6����������>�c(�-�C䓌R�[%l;�aE��UȜC9QX0���I3 �a���&H�bY�9�V0"BG�rW>%�������Nsk�
�_=!�[m{�{�����I\�r~`5 �d���W��W����~�<�к�0����ҋo<p���НС��G�wk��D��0����NX��[?��A�v��(kw[�������#�Fۓ��?f��$�o޴i${G�&�_
}�>G�|��2�3I��1I�f�ݖ�f�'�0=��wo����Ÿi ��M\77�\�mHK�V8IN�d�t߮o�n����>ʙ]�z��{x�7��y�5]�$]{	5����<�QX$�-R|E�\!Y��ƻQ~����w`�d@�,���
]B�������b�����0�e��/��_����.�t�|�+�Bg<'ǻ�6�TPj���;R�����e�[^VD-��I�g���	RD�a/��[�i~;>���X�u�!�3) `�x���Z6"��:�A��>��"3��_����*p�L��L7�_[��F��f{�9;P׻&��W��ٛ�+���?D����y�O~�O�$�@j���i>a�C�
rS���A�W�=F�p���M�M����jg�A6�v� ���b1�h��͂�[�d-W���*��U�w� ��a��P���P�,��\�+� ���XסC&�3J8��G4G�\��u&�+�S���:��t�/�[O}�Zv�_���	���U��E��!K��y|���{]84��,���`��s:FY���aK��e}kj1(��u`�􌈚����Pޭ�������Is��ReA<a�~��zb�G�v`W:���w��Q�kͩ�#S��P<��D9����d��'���7���Z]K�;���3�Ė���b���V�j���+{����c�"�[D[�Ŭ�`0?W7�/��L�=j�i�ℓd����\��޳���jg�C�X��U��,�Wʙ&g��V�T�(P��Fس�S8 �7��'�Q�KG���@FkA��2&A�r����c<J#J6@w/�5ޣ^���e糿����*���
�%9���5H�25q
*�h�b���V?y3��խ�H-�>[��T�.9o��9	���_F�瞵Q�_���w͌���9�o�S�eF��X�U�dc�E3�1���d;��}i!UO��)�'���ʫ,�tC�<�(�-��T�A��iH����V�aHo7�L�h6IA7B!z���x�-n�S��.Z�Ҁ����c�+Y t]����y�.��y,.�u_��<�y{}�p�g�I)�D��k&����D�X)ԥ�@с��H��ܻ��~?"	�"560B'���h<�׽�DX���Q[�AE����	&�Z�
��2�].#�} �v')��j(;����M��h?q�B/7��Q~A�ۜ��]#ٺm:��B�U<���D���D��a�V��4ݥ�8�7������������k_�BJ&�[y�y���E[�z�ʝ�YD�s����`ķ[o�7(`�1>-AVGt	Jg��R<��,u7��.���}Y��ا�����b��%�f�u�<)0Ll8�����>ݺ5�4n�0�O��������}����u�d�@�C�� �8D��>(�Ii9�����'�����9�~��T�4���������`ފ��������00ƞp6��^a�;#=:��W�t*?�B�yU�[�H�ʘ}
�m��Y5���S��SH��)����r���m�F��&2vIi������i����$�*��$=��I*��%M�!FW�����4�`��HŮ��I�
--���Y�u�y���_�U� ]�7N�A���#��`�w8����P�$����c�G%��Bv��w�	���n����>2P�N��^��u��7�(/�8e��k�3T�!�!�\����.�M�"� 	a�B��K�_|�� �Kי�����n$J�xK�>hֿL�p�ݐ����cP;2�nWT�ż�^e2<�׍r�x<l�z��Ǵ���n<^��q�{V�-k���7����S��}9��``�P�UW����ɹ��o��:Ox�`\Z��>@�(�����Nw����F����>�B�� 7D�+���z��-��[�&�f��OI��y$���C��C�A�A��A�5T$\�	�אW�pM��p��ƿ�:�1���F�!�<9�$��LjI���ι��(p��KaB@?�b��>r�RpM�e��Lkh�i�~���g{��"�78w��V4r�������]*_k6�sgc@�f�+l��㏪�P;����z؉a{��V<)H^iбU������X�E�ă+���FT�k�p�:��p�6A;�T��Ľ�����p�N�^�|F��ڪb�@mg0����'�~�AH��j���>~����R	>�¢���k��N�������@���6�gTn��F�$2{9B��h�ACy}t�5���6�i�>-<��p�K�-�w뷬%���\�FbME�	��Y���o��4Oy|f�h��g��;���+�E$8�n��?����Y��&�� `�^1!K��#��� nV�۩k�&"����p��X��]vɌ�s ��VP6�ȑ���}��gT^c[�E੠`��Z1t�|g�ӝ
��W���;�[��Ɯ�/�n]�I7\�i	��/��<�l�����nh��.p92�z�TW��l���g�oN���8m��ک!���:�[;H�,�:�����6�r��		���K�e�wӪ��jd������� L�� f���	���G�K��'�.��S
腈��cJ�nn��Q�U�t�
�y�$l�(��`���X[�X����׀@�oєm&��M��}��(!�\0�Y���&��F���bJ��$��h3��H\}�hNM XMQU��%<������MT$x��r-��]f&���W*��u��m\}��*ķ�E
Z��# MGa�IX�ԧ.к�2K�[�6S�c3���R�&�&��	߀p��K�sϼ�4gArj
�B*&/�47Je���{��s��ER򭼟r�p��en��ڪ�������+0#(5o�� ��+�W� �����sb�Zr�O��H��
�>R�5`�@G^^r,p����taw���>�f��W��ۥ�M�PJWqK{lp&A���;�v]+�b��p����n?{؛����iŚ��o�r����D.0�[��౻��+�!Eqf<p��6]'m��A51Go><!�*���+A�Q/��ώ�����5��W��=�7�����M�vo�M�\U��n�@K6���Dv��{�r!�Pw��\n��p�}T3J!?e+�]��<q�ph��ɧ)K�Q{� �C{Z��$�Z.�We��t�"y*=F�[�y����ЅN%�皋�u���*�QK	��S�`ABͪ��P� ��]�L�����d<V{�г}��mh��A��Ա��h���>��� �`���6[L*�lu8�Gl�[�JE4OkCeowqy#��0�6����O7��yP��d�����s�ݩ!WV�'�-NLh�h�饟���ի4}��(Ґe���%�t"�����C0F� �J~J6�AS��:�!bjĲh�$�)G�f�+�vu�Ѡ�x�P X�����:#ѻ�l��J�X�]^L�P���G#kK@A���{�����;>%�C���Ŋ1��2)�TE=���_���ێ�8��j8�h�T|ց`����O?��z�W��#~s!~v���=�u���{�h�;$���*�C����W��ۓ���]�b�fXK�}���}�؅'g��j`�fP����O<E�̵@��v����~���;����,��?3o렪QNO�	S$��r��%�+�p(�h��p$��O���4�ae8#A�K�����u�W/r�<�N}9�ϟg��dH�[�H���
��e�^'��0���F��=R1S��m*����[hN4�|�/4o�k�V�ѣ7֋S���t�WzI���D#���-S��Xq�ĔDՁ�;+I�a]{�m��P�b:���[�|���Uާ�N�,����R�cF|C��2�K"�R��z>t�7�	͘��@_8S��#1��v�����C�ߢY?}��w%v,pN0?=acА=K0$Tf���C�k��鉄:s�BI^�^�I�W؞]&nR�v�-�ECY��lM�ǭ�VG\���cjGhv��'T� �H���a�G=�����(̬�>kd�b�Ѣ,�qϵ*<Gm:Љ,4+,M��/aTej,d�S8�|ڟ�)u4m �:���/��c#�n�2g���$"����W����_�7��cr���,�)�x��Wq�{k/bv��2��g�ˤs_QV����x~��z�hU8Jq'7�eq[�I�pI�B�����_ʆ+vkl]��n�zr���A��7���MRS(Ke�L�^\ʧ[@�����������-jߥ��Ւ�K��Wӂ<u���TH�$wI?�ӯa��-XW��ç/�ӹ2x2C��Сp?�������>w���S���PZ�R	�r��2����c�9��G��Q�
y ����O���=�`\�=H�������E�]�SL���3j$�J�?1'")�S�������`��lH�5�Ѡ��9�V�c���ML9!C��#Xd:����=CedF�1���k��A"hl#Ho7U1��v�pP坍�־�������!��,��}��P��,[�G<AC }4ohF�\�P�tv�c�ub�=�"��*Q��NWA+�V��n�#'�̻%¸�!@P��z�u��~"0��*�b�J�u��&�t÷��.�j�"]�#Ɔe��_��-���#˝��,�7<��1� �t}g��3?u�3�YlR���V�ps%���ǟ��U�:n�*�ɽ�4Q�@1.���;����6���
~Ke��˳'h��q��x7A̐U��IE&�)�ݚ���U`���)���
�ܠ�lx��/9a*e���Q���\�vF�y�Q�"R���Zq�IJ4��P�&>�H����:8RȰ��E4Zm�w�!"e�$�='���B�9	K��r���V
�5��;9CV$�ξ�4Y�7���[H��7�����pcᏒ�^܃���F��oFq�	����/��u�aIX~�:G�~�8�<y>��hs��=+՟�X�]c~�@7O�c��+� �i��Vs�*��%$w��S���,փ#�,7M'��遃��!gZ9Avdi,�E���ʿ��7U��!�����@�Ne�fj�3�L�5�*�ֽ ���a�T��1f���*��Ƃ��>����W�{,�WQ��F9o٨b�� bL�3yc�X�
��f�e����6z���,�G�/E��f<��&�6P:���ք8�W�\~��)���wN`�b6U>eE�S�C��7 v}�1�z0�"�� �X���~�:C`��38�$�䆔6��ǆ��=\\�R$�_h@���r��n�U��a�c=��U�x�u�{�bD8�j%:�l;cg�\57K�G(���%���]�w��F&�jz�C޺��r������y ����6�;k��R���|���
��VJ�[EUS6�OIzl� Ԇ��w]��Aj`����p�z	�G�A��|��x	)��څxO���Y��cX-�K��"^>�#(��M^m��!�� ���SCfǮ�t��2���A�j�J���'����k:PT�+X�!Ų�C<lSi�i�8�r���?g0���w�����v�L�~WX�T+����Cs�������t�����KL�O�
$ܵn�G7�e�y�Paei�r8���x��;4ɩO���j4m<�_li[θ(��u�c��]3����2DY�PS�R�N�.�e$�;Iz��;�>�f��{��_ �����ɝ��d�B���3���|�B�ޟ��{�ݿ��҇��zm�����;I f@!�4+���{@Zq'Z'�T��j�oO+/f��Nz���%-GA�xc�"�7��w翬�$Ŝ����A��ຂ�QH���愡�{�7]���#��������=qĕ��1� �z��9�g���L.���1��h \�ֿ8f���p!�����'U'��_�}cU��� S��A�;��j�����Iw��e�ţ�6vY�BK�H1{�`�_�d�W5Ӭ�ȗʄ�R|ĸ��$z������H�.ǟ����>T�{���ւ1Űd��%�c.�Y�\�c�P7�8&�Wp��DjȣH�S�n�`�sP
I�����<��� o=˥�j3��E����[������`�7��7�t;p�/l?;��&,9��Yd G��Y1�3NPQI�D̃D�e,)�ܲ�>r�sLu��x�Y����%�KtQ0 �ݙfY��A'�d��,�2��k�?VOa�M�d�ي�Q�c͎��KA49�;���Jė�B�[I���1rw���S�TuJ-�*�)�*�b��q3B��\զy}Է<�M<mL���[5;f��7�ߝFd8���iɨ�6�U�K���OQ�V>Vv�`0u�ߕ�v���vWæ����U]j"����@�@�n��W�m���p���f\��7�V��Ԙ��G�PQ,9.U��T��;�0"3^
0�+HS������˨I��(��S-/�������7�x�{�w]�!_����V��$���Bˑ0DWl�����E���.��S8v7�\Ճ�%�
���CؚQ�������,��b�@���;i��=�,�*P�a�6# Q�"a��B��K{��s�9��1?I0���Uא�O����/�F3��ȨI:Z�@f%֤@�m������ltgY�D�*����'1ͳ�$mc�a^~�K�IKpUi����Ji�qe��F�"LMB݄G���f�b��E��]�9*<�	���N�b��0xp��y��96�����R�}O�!�oBWl]����ݑ��T���q��m�M4�Lb6׽Cj,��B��'�p�������y汊�n�q���Qd�I�����e�u"��m�.����e�W�ҿ�qX��X���ސ??lB���o<�{�1�r�ry^-X��ǋxX�;5=�[�2��o�m�K�?�̔�,7A:����ԫ,����D����`+A�ԧ+"7!ܷ%�#`8?"��\c��G���R��<��5f��cJ�ٗQ>�v���D�z�@����Us��7Ｗ'_܂/�Z�p��Yl!"e�xӄ� ��5��\ǟ�Ns��ir��؉��k(@08�د��맙����)����ΐ�����?#oOC�FYk>.�ǉس�}��\����h�v�{2=;n�6�\	�|�Z�s!�L���=�́z[�n����0ꀢl�Z%�����+�X+D�����Z����P}�o1*����n���M�֋�=���7T*�a_p�۬n����`[�E%/hҜH����DR�y��z2b���D�@5�*EFuh���Ј �Ǝ�a�}��E���-� ��}yNk y&;�	��9ڭ�D���;���R'�Q)�L��_E3�� �_k�Yp�=��6!�a�4�e�;�K���u�5z�B߹	{n�2K.��,p�e<�gNg.ӎ�'�(=�`{���/"����s\�N�����m"O��A0>�`�vLƗD�'�My���#���o���n��x5��o�-���h(�?���jY�z'�Wf��Q<��Id>@�ϗ. 5t�c�'uN5#��0�*=�"�/dgt�vO���B�E�z<��ů��?�ku/ժ��i���j�K�i	:��y����}����=>��\@G���E��kX�����uzC����~�zZ�4!�9��(cr����s���_ ���M�to�[���P�;~��d��R�(y[Kȥ�N��T��9_��c�/�4��5��ӧB끤a���p؈��v�!(�����UHڮs(���&(Ǥ��ni��KX�
�9E1����Q��=��4�m@oPJ	��j��"Ñ�ߙj}�B{1*�W�j�b�,�I.ݒԗM��PB�=9JD��J�	��T&Z��x�vI�L@ܢ����.,!��Q��q�ru�8���61���8i��Iag�
���SHGYO�0�[�k���Mo�����ǳr:*6/�Sī���(IܫeCK��2g�*έ�B����wK����?�Fq6���-?U��L�0�(*�!mQN�+;�)c��a��d����l����%�i�N��@���#�&�b�rE��|}����ؘ?�t�Rǅ.U���_�2p�`�%���v�3A��l_�N�p8�]2�|cy�_���1���\#�b���8���KnD�hDG����h�S_�7 g�|���+�K��+��a�7-KA�X�`�$�&�D�&u���!���Y������شY<���	c� �t��<~�z��w����z��|�c\�P�TUuzp�y�ș[��h�K.6
Is����#ʦɰy>v����|���Ri���o�%g��}ۈ�gy9�K���MYƋe���noboH�M���M�l�]����d��	��e￘�o�����H妣���E�������2̅���� ��h��?��u�ɘ��1�Z,�kG�~ֆD�R8��De����}�G8k� L*F�J���l�Գ�V��� �nGCb�u�2�J�Ԛ����3�y@*�+�2(@e��-�9�ӎ��Qko�����3BڲRF<ŕ�P�_��ª��������W pd�n�l�"�͙�Q�I�(ٻ�½P�r���ىW�C���6�@��.0��>cAU�V�aJ�\�àr+����$�\}� �̎ʤ���w��Vy6�2�I�M�'�����I_���x�t�K	�˩9����7��X���hfʛ*��u��7�f���x(d�XJ���f�����~1�r~���F	�J�s_d����Z.�	D�i�8�.r��عq�&�-��ߞ�IQ�1�ێ��p��:�P��P�L3V�e��M�e1U-��+2V��Ԩx,�ȥ-z����ğAԹ;V"Qpo�d��a�΢;�|�Ҹ���D`�:��Nw��#$Ӊw�\�h2�
lR�t�D.Ì>1"V%<�;,t��Hr��A(�x�A��t�]4�{�V'�9�̭��R�}-u���@�w��5#�7�3�{ �1�"sZ) ��B+��@� >�Um�w�\1s��>)���1q�����B9�� !`�:����Ҳf/
�ME��֢�;�L�H�#��_GQ�:��;��Ɗ�ާ����Ԯf(� � ��Dx�]�(ڱ�3ǬA���vt�Q�ڙ�SN_��ә́&R���>���O�_���<�;�wL��V(]UI��4C\�����;U��da`�H���OUT7$ҝxf	�ky��?2�6/LF�i)>'��LE(g���.���Ie�*���~�f��'CV�t��4���i��T�0=��E�T��OUwV& ۅ��ܧ��k�ҝ���)2�D���S�s8$�����Ip}�OwM�M����xJ�F�����C5k������BEq���m���WtM���.�9ȷ�`/P`(���*ω�,i��M��MW��C�9AA�4�gH�ģ4R���8KI�s�!���9D�@M�`Q#u2���kf�*N�8���\�Ϙg���u�5����kF�W�R�?��ZI�0'��g����Qs�-����>��\F7�{�αw��za�,ak޸�`�愂��"�G���~9�!S
^�Dk��qP�5��ڼ�ކ~���_W�62)א#�H'4)�+�ky�	WZ:-8u{�C)q�A����9����$�4�ZYIt ���}s-t�~K�lֻ.��'y�Kh�S{'ǸävG��B���U�1����`ʔ��0 ��T������0Û��|�Y��礘���wl���A��X��,�&�7��yx���6���9���&�|�J�m'���e��2��

��$O�����f�����D!�)E���6��;q��^��p�_v�t>�\����ϯ�a�M ��\CR Z(�DF2/zj��BS�l`�Ȟͨ���G�r��OX�F&���;Өt0���:K�|((;�9�Dypc�%ae�fUƥ^��%�$���g;e۞yЗI�V��N�5��6������5uL�vr.x�,���*���u��^���b�?�۽rkp�#����˫����f�G߫+p W��c��֟G���i���_�J�y��S5w<]r
j�� �|@B�	�e��4��
��B��d8��!�/&�/�1� ���*��ǂ��
��2��Z��6�@kW��̽�ɂ��/)��u���?O^C�K��:�i�R�����;�>�o:�Ӫ�q�����s&�'Ѓ�������2�ǻ���e1�O�ĝp%i�2�i�W���~ �b/0�E]�ܜ�8JYL_S�]0�PG|t]����Qz}�`@�+�px�'Չp�`j~���O�&g�����[�F��jz߾�������uU�GRE ��a�eRM=E�QCdsF�CTa>��j�������S����>��_��Բ�Gt�f�	�%j�R.�� I͝.�����8y!�Y����q�8�d|Jd�\�*�Td7�&���������Q91X��Y�[�Uo��p�־~����>���{2�������*��-�Է�P~��4�{N���t�
@�+��fO.�E�����Ȕ�mSa3Lc�=M�|�μ�˵ЕNz�X#��Q���5���YZNR�\ �hh�ϗ	=�ʨ�����g?��]Rf��cI[��O��h�Ǻvq@f���\�dX�ߢ�� Y˳�M��(��U�#�F��6�b$\�uW���-��@
���?���\L)�1�N����y֜H�e�����>�9$6,%�y��@�gҺ� ��7FP�2 %��
l�t�=-<�^�LE��x)#ن��A�L�nby/�d@�WdC/eC �ɇ��/6�m� �M���Pgk[5��uW�^�� ����Q�p?�)A�+hè��5�-xֲq����ɶ��J�Vn2��W�N%80�`u�	�����7q�#��E'������ގ�Sl�A����_���Pò�����&�P�@-���Տ��(�Sx�]��h�����X#�b����s�� 8�@�A�g�zۡZ�8��(��!�ܭQ�\�Y�C騲�j_�x�S/�L�9h4I���yp-� z\��NoT6�������x�%s2��	������c����VI�����ۙ��xq�a���S>1N�\��{�~�`��i�(�Ϙ����2�?����w�T��GK�k�!Š{%OFvv&N��;�h�� ��Y˺����gxNlÙ���>h��=�T*�=[�Kb;	/�M�RIEMF���[H'Wlj�G����%YfNY�Y��)Je�=������؟��پS9ۂ�蘝z[��3��zHDy��n���hʎ�����=�*�0ԋvo%���_4���x����Ի��_z��2���R�ݖ'�
�DN(���p-�t�<˚��SxK[�q/�0��)kw�����)p�s@oy��S_��_�[.���~i�n��;PI9xND�����k���<��c+�@��U�s���0p�QX^Yݘ�f�#��KjM����H�|��4�M_��<��W�8�̢3�J o�`ǻOnT��?�i�:*��\����-�X�,��L���U���>x��°EQ�����rG$-��B?X�A�"3�.���\��7s܈���<������p��8�6��Z*�)��A�v��ڇ8�k��R��g�e �\Js�.o�pxϝ�#�ӧ����u>��	�v2��#DRg�t����$.٧�}?�2����=!Yx���%������_��e=Y��8�K�fS-��`L�0�V6���
��`U�抚����ܱڪ��UA�����w6v흽d{H���;�0�����ʇW{��� �#���S��:�q|�RJ�L=���ܖ��B��ڍ�MO�F�9^=��j> 4�1L�Z9�_h�s�wp�H�ҭc��w�V�|U4h�����Q�����U�cM����Bc0Y�ܾ=|ݠ���Z����
Hh��[��	�٤{Tyqqv���C^�7��p��38��emՍ��,���$
� (^���P�o��~�9��Wg�MSK(�V��v鐠yT�gu��Yb}}`/}���;Dv�D�vJ����ط���X2��4**�Tɲ��
��{L�����aD�$��|;��ԁ�R�N.�lo�lw�c+�Løs
Ii�C9ISb���Vhѐ[�Au.�P����˔�?�qK}�?+s!ț^O�"[g#�d7�Ч8E<��[g��������=���"ٿ�i"0)���]�U_'�Г7e��g�L��S��Z4'+IT[�f�(^P��9<��(2S���n�j:�P2�2�[��W�1c�΄I)�F(�*���O���z����V�Xl@�?@����`S�ϥ]�),��8֤F֬��h��#�rl�ƍ]�?ϒr�Q�Ś��7�e�̉N}�^gU�-�f4S�ߏ�jm��MT����y��1�f�wf����~�K��r��4K:��D��%��%�l����dHny�
��,r
���)w�ߩ���un�tLW���Q�R��Zar:8�흤
�Xr%�dX�pz�biF7=x���v!9���n����&��o��U6��ð��K����&}���2PbdԿT��#��N��u(��޼˓yU�B�Y»A�_X�&$�c����[Q��OV�R=���N3��8s5����9�tF3�|�56�"��Ϸ�u��}*��С'&k�h�m�V�$���pSY��mN�hNq1�5�M1�@J�� ��A��T��n=z�H�Ik��qGS�:O�M�}ir�tY���C�3����rѠΡD��t�|ґl�a��fĤ6�Z-�Hћ=K��dYS;~:si���E@#-�?\��dy��e>���e����D�P�#6�r��
�v��a]м'�5գ��͉U
!7�� }!. ��:3��m^֙]�0�9�R��f]
%�}��20+���� d,L5��VFܲ�EIž� l+���$tJhKA%�ݰ'y8I��5�}���ʂi����5�m�T��U
�ƨ�@�Hua����I̢a�h�C�ց,���D�~�4g�2'}�k�4>l�#���
������Py72^(yn�DMs���!�������»"}�iaɖW�GqR$ٕ���¦�0Yd�9ƕә�,���#{���4R��`5�u�(F����F*�_>�䈾9�{�w��#��gHݮ�?e[Vm���kXf��ZE� ����M@���9?,21������AA����g�װS��]�_<�v?Ƞ�6�ۨ;���n6HT�?�١���"(�����}����_�	4��B����%�ˑ��S����U_���3��K�>����[�Wc�3HtH�^ާ��Srġ~��+rg�X�ZU���Ǵ;�*�������=��wx�b9���F1�-��� �ѿ;��T�ӓ��j�^�KBԐne!��;�cd���^l�qC)��L�I0�NR[����V��q( UB2�/�A�����LQ��T���5;�W�@�"8�&�<()����eg�1m��a����1Va�E =0�5[��#*
[���潴{"c�}ӱ'�ˤz���LM�[#�/��a�&M��~�r���5���2�BG����/�)���e��X.����m	SGp�T�Z�x�T����f���LZE��{З�e'%l<�~���]��������Pk�Qv|gg|������%'OW����❤h3��U�0�W��a���p�,�cfC��dwR�	�1��8Ȧϊ�($���m�&
�ۘ6�����~:�Î���/�;����,X�:o@���Sb���<>�Qj֫6m��}��j:T5��,n\p�g՝�}��p��Hy��k�6��3�����ThL����7
���*�8�l���Ra��/���7w_��!!�U���o7ͅlu
�E���#�Ω�3�����\�	��R��G��Sw����!��ڏ�4\�ɇ����fl�c~��6��'WQ+�Q��!�:��6%�y�l@���*���ق,�IFM���d����1�'�rvb{�r9�ә����-(��eޜ��p�J�B�5��P�|����s�LQ9�cg�1�����z@�~R��u�[�ݳ��&�JUs��2o�Sw%
G�n�
(BWSw�8~��G��i��؂΄��BE����+�I�j�+62N��B�%*a�uC#C�v����\ƞoPR�	�0[�ց��[�4	q����V�\��D���JR_��;�0�T�l��f�(�}0��XM%�A찇rr�[��5����)�z��_NLsf��zq�8���^q4��ŧ�#��/(5e���	ދM=Q�O��h-.���"��C�9X�<K�E�#�/D&c�>���2�:F�Ȳ����-!>tAb��+�S�Y <�ۑ��l��]"�!tRC�ڰ�v�,u�m��J�����~�4�ޚ+jY@�fv��0��Vϧa�-n��_,� �0Kc�m~`Q�aH S�p07�W'ާ��܇��[���{xA��.ܮ��M���cq�6jdp���۹�/L�k��T�۫��db�	��:]��,B)��^-��q�S����+�X�.�T��L���I�=���D�k���G���WN�z�@�����ɑh�w��-�^�A����^q��&�@2��n��iIܪ��<5���k��O޼J�r�e������8 7,�8������2)<L���oۉ^T �X�jIA	Fz^��_��@�������0���m�f��́�����eE{Ԑ�x�ޒ#��q�2Rn�dkėo���ٍ���M�0���z��C4D���GI4���mT�緧ؙ�O>�g�J�L�V�������] �VV+t.���}��<�
Y��\_JAXj��fD��ʿI���jڥKu�-��<���H�q����NX��<P X��?��i{������y�)! ����̍�\8C�Qf��$1���L��{*��ŗʤw�k8�#T�$uT|�{�$�C0��m��1�Q�ros�/G�-w���q7aR�	��Xa���6Ǌ�+\�$�����R����˺�������k�G7�<^@p;�|cJHn�ȋ���t�Z-��HgJ�ع'C�5�P���oCG�8�)K�����0��I$.��߃��3is1�:�*`��Y���Zt��8�4i}f2gP �F*��D;:�x_�����(?-vpОKo��*��̢<�v�F��`�`�y�����$Hi�X�e7)�*Đ��x�]��X }�8�r44��W�qCi��5�2��<(b�8�5� $�Q1�#+~Ma/�XX���;�lJ/�{Mʨ����C�5a���O"�w?=|���y㘜�6x��r�����W�s�Ԉf�$��T���>g��I�5,��J~O����gr22S���8�@N��Z>tV7�Y�)!�����T珇@!�2���1�͆�a�g�!("r-��Ճ�-��%���p��!�\{<-��(!�ǈ��͊�]�|�R�4��-��V:#ֻ��B=�=Y��x����Hx�|%��Q�zi���0S�\��~u�c�ra�x���s7I��1`�f�tJ�#�Zk2~����W^.E7`=�T籎����C"xՋr���DY���6�'�Vo��0fSW�g��
��wͩ�0�#�7�t.MM�S���-�s�t�Wn�fe�}@�!�4� �v�:s����[�U5%���8�C�;�e�4#�r� �X9��o
�9� ]5�_mi������B���wJ�}= �d,-ȗU�ŕ=��0���c-�5�t=8�����Oa@�
�����B�RfE�K�w��j����Je01�J������b]|�ܧ���bp5d�J�:��?(rD�&�|��#�W9[�iN5��mǛ!H�U�2�{��N�/�4�ޓ¯���r*l]�?G�2ת>d�s�ͩ�cB���wa#v݄�E����v�Hj�ٵ�>���?��s��n��R�I�( ����;ź��E�[��2i���iػ�G�'?ߚЊ��3c�~8��%��R�v��^x��� �0�{QF���<`��^a~-DmC|�M�P��]��_i˵�N�;��b�"���k�ڀH[X���/�H��_��D	�ЛG][�*؝,c�p�TaLf�>[�.���Q8���\�a��.����?�z��K�5��D�Mrx�s�6w�N�1j�*��_G���4�w��E3�����/G	�r�٣�H�}�+�����;)Q�B��^�P��oČ�T����!��n���W	�?�EZN�wF�k_9��5�u'��Q7H���{�h����I��Wܔ�bL/���̧I�=}���6y��t�N N҄3e�}�q@�
�"Wˬ�ס�N��}�+�U�dU����#���y?"��d9����Đ�I�3��z���2��v
���,D��|�y
�R��(�X}�7-�?�8�������}�/~� 
}��"Ƽ\8���כ!A�@^���e�����]�];�j�u&���DI0G�Jl���_�D����>^���fϳ
�����+^��M���%�Æ�m!,�ndu�ow`Hqn��Q�&i	��#=��Ǧї��0�����x�� I��	��� ���s:�n�9����%!���q0?>W��=9�9����Z-�����ȼq�1���j�*���C���	V؇y���o�6[�V�,�A���G��:H��|~C�����+����'�-�ˮ�?��@������[���I=s\�gOqf��[�S���n�G
���%�3�_�9I�oz�"��qg���n?�3��j,�F3�`<�'�Ru�o>�U'*%���*P����Z�����~��;!�зxF�m�Zw�C��2{\jq��]��T�IZ�Z;CFV���I��)����蠤�Q�)��E)���:^H~�LA9͚	��!y�-�A�';�G�%f�y4�dS�����Պ�-��:�jˢ�S��~����\����jv��i"�r^���n
&Sl�HG�z����N�pt� ��<i)W �$\v�-�<�gu�:^����X�<�G��<�%�#gh���z�к ����nd��ȹ��;HLA�v#�Z�o�芕�����q��v1a�M|��ޞA����c�Ff^RT��@J8řwǷ����N�ySʛ��a�;�{->�j��=�*��/)�Y}>��>���ꦰD��T��5��;�TX��[�؀8�
��8W> 9��3����u�ڼ!�d7��55 'jh���]��᭛�(N�y�=�FL�i+��8i�v�fd�����N�Tx���A₋��ͨtg�{��#EZB�|ɇ̤AO `��'f�WM���Ca8G�2�����wN+������Zd=�ٹ.�4�6�d�����T��a�c.��)��Б�=��K �6����v汎��^HE�^_`�w]��\)����著,n���sf�H0YH�!]۰V~ů��=1�6���2��ĪXgA�V��7�uQq�7s1VY�w�H`�D�8��4G��n�lg{W��;a����bz�X�s�m̖A�L�6��3�!�C,���x+�i-�I���|`�|��{N�0b����͘a��e\��i�y�iA&zL�'���T�2]ݴ��7%B&��&K���?��
�g�9dH�D�I�<�_:��T9x�� k��������!O}�[0^�Z\WB��i��0�X*��Q+�����	tEP�P��c�J}0�
|M��;��.�Ţ=���@� ����x�a���_hp�W��Ľ/�4,�K�kq�V��S�zj�X���nTb_@҂$��$�p�Qݷ!w@���r�N���`�Q�f�KMZ��w��$A->,�X$H>�]�ҵ�D��:s��*��1��JC"�x�����N-�My_aX@g��/�sK@�"������>\^�^q���*��a�&m_�z�-�z(�;U6�c�g��f*��q��e��}�# J�Jz@a�p!��	�#���6����)���=����0�&^=�q���~ɨ�o������cu��xNž�7�Ǥ���Q�[y}ݿ�����tޡE
H0i�����|*���x�b"�g����?q܈q[��je�ѭ��C���3��4|��Y�b{�ʇ�"����2���N�RG9�w�";%�ƕvM�u�3���<]�cor���B6;�37�.%���U4�eH���	ިϨrȪ�u�5j}.�����kpsS�����Z(����m�1�U�\�TWehd��Y&8�d�����?�[�=���40?T�R���n	sfu��� XOj��=��(x�G6E���0J�C�P�h�޹؇&�~�$e��A�~��B��Rh��U�	 �d}��b�1H�%ESd��蝥*	6j�Do�C}]e[޸��°��2i���J���Nּ;ŝT�Q�z���*���T��W2�L��-^R�b�81A-�l����p���[��}�X��S��-���6�Scxj����ء`\�`���ڦRG��B
�v�H�9��ݖ,v�����C܅�B��P���O0�����t CAK���Y���b���ݎY7�""f_m���v'�-�Io�r�:,�~s5mE-�G7��t��U@Z�:���n��ֶ���۟�d�'�닳�F�Gn)��т�����&��<�oKH�qt�\p��$��צ��
c�˩��@GxO�a6`�.���tm��f���c�?4�k�Ru�@İ�5�t��O��|Ĳ,����N�4	�@����t�y"��G�z8H��b���w�t�y�4x"��1�o��2�/�t� Vǔ� DG����� D0ؘ������Z`�;����c?�?��\ɷ�2�����W��?�x�~��#��.zp�ȬZ��5JѰO���³����3^ʓn*�2U�?���V�|���݁���n%Q��l&Vf@mz1"\�|5ɤ�C��P@�W��YB���z��&L*IU�$��'��.Um���7��[�R�`���9��ʷ��H�>�JOz����� ��`v�{���׳O����^����JN�CvSpi�$;XAJ�m�L��z�CU�u�6�\�.�C�͞
�	���G����T��V�rV���{:���{�F�h�f����Xu�I��� ���h����x8�%����'��n�K'h���mEHݏ�����Ȱb@f�~��M�:��W�/�e�^�'����j~���%Ӎ����%��@7)�N�8ӴWl�r���_��e����S�عßݛz����`A��Krb��x����M����i� Ì��t�|�w�v�A8��'�!{I���Q]�c~t�*m 6���@�T\Qc���#Pqӄvf���α��kq �\�xͿ6@�����J���֗}����
�xҍ��#ҺY��~E=Mt�濪7e!����C
�?4�l=<o$�0"�����g��c�vy=c�0b}Yv�(�5$�U���R��^g|��3JZP������!|�"\FL�9��%���R�J"�	�U/C�;	
FE����P1߭�.�i�A�����ئ��H�	*h������e�p��$�S�#4Z��RQ���9��g�ڸ�B!�'-��!
�D{[�xU�KpB�$�SA���k��5ݳ������Y�L�ҧ?2��P���X��Q��R�)�4;P�U�(d.*��x�K�՝�i�}D�H�.B	;U�vqX%���~��e�z �;���	��, ���j.�J �����g��q�)҈��+_�$�x�ػ��EdL���h-NN��T��t����$��Ͷ~�� A]cP(EL�A�5����MD;-�MH��eH�Ā��TA�O�W�L�s�E�Sg�;!w�	�@7�H��dA���������	U�@�h�=���?�L��I	��q���OS5H7Խ{ �IE�3�"'b���'4
[R��Q@0��r�f8��k��@[Rr娲(�i�!l�^��p♇߶;����^+�����q�U��=�����rX3c�f�x!�E)���("mEZK�I[��P\z{����}�p�˚�3J���Z�g(����m9i���%܊h��5��Y_�Y�_6����;��
��|J	)��;m��
.#(D)��X�n����4�`�����?�ԕC�Y�N�o���4=�3����c�r��.�*�L51��<])A�C���sIo'��^D�T���1���
+�Ώ�=�B�(Ih����N}1\�B*A&�	X�e�]����,�G~]W��,&jݛX�n�t�a�������8�z����-xK�n=����P)YPe\G`�v�>����y�B��z���}O;i.��
ٌ�7~&�%%�c%6M�����2�U�F����+,Y���@i7قnI7�rMRՌ^<44=ICzs��
�={7�s���,�/k��QI��-zg�R�
u40���Jo�C"��m�����Y�"%��F`�:��/�=U��j�tű�O�F�5��f�d�4xLV+t7n�N�op���O�P��=��I�&�j(���m�$E�jS���d�D�@�#�(�ʹfb�<w�c�%+��c�X5+��W�Q:4��Ј ��hi��4�`?/ �I���N��)5���4��d�~�^��ec%�ࡈ%�T�pg��ZΞy2��*(pn+yY�ç��k� ������5��4!�<�1�'v�]��:]����1�F�1��1����u�{�k��yb9N���������n� ��d�le���E�G��(
��m�k�"� �9�Rj�ӥR_]�l�F�F�)}��BDVY��Ɋ��j��M��D�:75����� :��e��l �o�RQE����6�BS��:*��l��i;~��ti��jC��N��8"���K:|/AX��d��f��Q]�)']��I�����d"vk!�\�3����P�F�s��Cn��6��:T�'1 XDŧ���8I��K2 �č��^i]������Tb���:|���P�ɓ��'�ʚ�Ο'9���F\���/-:��
�����0�QCR�iD>�;��?��$n��US`+��l*Ej�W;�)Z���,K�XNs�3홃�e����jf��c[p�d4�^mW�fZ��E�}ӈ��o��"y�Z��3Dܒ,�̂)�E΂���T�����]�c��=�V�LO�dխ3�4j��k���z�V7-�:OxE�n�F����d0���+e�TB?����b���j�>��;Ez�j���1Ц�S���F�{k�]R�1 h�����KMT�WS�}���mM��/ܫ�{��]�Q(>E�T�_�ܤ�y������[��sN�ܫ)`�_�e��s4|ɖG��4�jܣ���*�J��fǫ��0�(H5&w�����/�t���+!��Oa�{K��q�2��rn�׷�a��ꯐ�u�~�*��+��i2�6C�7p�@��~]�G@:zHf l%5�0|�a�Ţ�:�P�������6_����F��*�E,�l���[�7��޿Z����ܒ�H,�S��>L�r�o$^�����-�L?�����IFȫ ��[<;Q������w�Z�v���C�	Z�W@�t�N�i��Ѫ���`�x\9�Y>0���	��9�n���������4U�BU>P��@�l��Yy.M�+����*��
ga+y��� ��9��lp�"n�z.�O`jh�M>����`W�&^W�"����ӻ'BBϼ-@c�0j�^��
j.�AN�=i	#�l��Pb������51	V��d(ɋ,��V��bG/>K���@B���m�?��y/Cu�h.��Mt-nO���f���#}�z�)ڧꥌ�
�x��O���O�S��3)j�hW47q<�ߢ����d��������Ϣ� ���!J�q�A9J�@v�@rͣ�ɫ��>�a������-�r�}չ������k˶��i�!����c(q\�b ��ua$��C5^�y�ۍR]��������Ä�<��W�9+��=�ON�C���I ��u@8kzB���k9�������߼��&�����Aa�i���"Q��崨8I|��Sl;���8Oԓ24|\a��&9��:�8ڶ`F�Kۖ�N��m���Z����R�֫��{6] ^��>�l3�`F��X_M�vV�����C�)z��1�l|X�Ť@�/+�*��t�W�W� �eq �i�#��'}2��:��Am��uRB
F͋߅az�� � �:����j>
y�{8�?�:"8����~�>��TW�XŬ�;�<I����g�
mݠ|�+�N�A�|�*^���q4�M��Gl"�K��$�'��?#ᧇ�ȥ��h,�u�[���I:����S�;�_O`�/�9�k5�k��P������+'�P��-�f�A8C�>z��n��n	D�/L��k'���-��n�x�*���8��w~���_�^�@���#:2EFUϞk��A��M8���3��@tm�vw�ݧ1�=��ܼ���؄�4[A��EEHtV���p^#��e�Z%m�n�{T��/��@�Ӱ�)ș�l�[�Xo+Ӌ! .�!��9.�®�b�99B�z�B�
���tjm��
���V�K��{����b�}�F%����w���Óaճ��V�����9e�NbKF5}~���/;�]jl�Oe���֭�-��o�G|��J�q:��7'NwrUS(.�K�I^ʚoʰ�G��5�4���=
_&�M@;��vM�li{*u�?�Dbd��;Ͳ�FڸQ�P��)͙H��� �H*����}Dr_N�,N��cT�^��wJ�	6���[��2}��HB�ɦ��᧭l,~VAF&�MڴR�ą�^�ԜS��)	�e��b��'S�u��ޅ�+<��b��m)�����ҔݘT[���0��e�P��Z��&D�{���s��$��x`]��+~�K8(��B�������G�M7�At��l�\��Vq�t�1�r�UQ��\���.W�zٯ7Z�E6) �a��^h����-�ԇ�1_�.C"��h{ݏ���Z��/���{�Dn�����9����|N94`��ޗ�/p������1ѕ�nw��ݿ�)��])��TW�Z�;A�(�n��/��Hm]�8c�_�~L�z�`O��E�3"�HGu�T�q�'�D�U����1�S����j�?#�,@F<��o�%G#]%"-���Y��q�l���~γ�����7Z����B����� R����w�i��F�O�����.�:KLi�81���5��@6�,�����j�xZ�,���=�jT�(�]-#�%`5,�[��6��-��'ۓŅ��jQ��L�����j5М����Ƕ \���3Ż��l��办Q7��t�  Ů�i�ƏLCN�[��q�"�6��0NGx]�0�Z�X���tøxS���f����2���T�mfT��Şn������UqT�LJcr���3��PH]%����t�խpݗ�_P"��cx���� J����-�&��M
��������`���%�.�J�!��w�*>b/�F�L'Xm�:��P��w�'�a�ȭp�A��]1�����C\
�3~���^�54�-��_!�I�Z=T���n>)�C��c6�i���8���4�8��f״��7�vM��E�k��>$c�yz;K�؄��.��Vi���M��!4��j��d�_�]q��Q>����wp乨[�%J�z�U����9�x��R���	��=T|*���@�`�'�^ ��N7PPF��.��DO���"w�n<3Njw^�jMq˱ss^�}���z6a��UVou�pw �0�OK̃��.7����B%,(1:<�����F�(;�����E��	��x�i�/[���^�ȯv3kD���&�T`�S�$���A�A��������˶,�:rb�so�����쪴Q��j!{
�p 2�쳯�d�Tj8�!w�G@��ڹ�� �q����d�0��IC��C(��s#b^	�Ī� �]��7�&�6���2�Y��Ġ¨N��<�p��d�)]EJ���� �i��ޒ�@q��
���7j�:K�0�kb�Gy�:V����y\��
���`�XY$���Dh?�i ��g��/$���x/?r�b#�^� "�'���p6p�``BaI�Ra�Ѽ�;�h#��l��-@q��q�U�*��*�I֐wi�t2�t�}��8X��~�F�ּ��P
�6��h���"�E��N΍���ə����(?4�0��]c:l���]��ƌJ�҂:Aʳ���ςᲜ	9�	��[a�����;�Q!%(_ˊ"�Z��E�͵�z�XF>���,ro|x  �����S-am�t4��nЂp�����P�O'��s����Q�d��[X��fq�SUb�$��̺ :�=��<�nw|6�NgSϹw�q�
�ky��x�?p���2�c�mg�O6t�F~2;���T��L�������;��W*ޑ�Yn�Q&��^O�e`x��M LD@�_���TstY�g �α+Ay��[��Qh�|�T�5�e	��h��O�z��.b]�CWv�|��"������s����ܑ�L(���af.C ���_�Y�8��E���i���B�s�*���K�(�Q�L�uq���̤*=�Y[Uou�� ��lc���.~��${�p��Ճ"�B��	�[�>mͿAt�	��L5��O�Zэ�S�@�a~�ߚ��a�l2��=y�S� Ҵe�����ҍ��S����Řq٠Ia��]�� [b�+�B��T��:0\�垟�Z��]'�}ڹxU�?��S�`��c��v��B$��{���+O�qt��B���&ƈ�EmN��6���6��t�v�0^3�{x}>v1|��'����V�C�fB�p�v��̂=-�R%�$.�S�޷�,;�/�q���[Ay�}����הA�:��R�����4e՗.���Y!b9I��jH}�t�fIeI�"�IY��2@���^�-�'/K`�͐S�ǹ<�	�׆
.��YC{�R�JC��t/�2�M8��'0��x��aq}��i���:�&��Ed����+��v�a�0���}�P9��$M����pV�6-�e'��U+4��e�����������b��Ȫ���)�8��|c�״ n'�M+�f����o�(�"
��� �⾼�1�:�����)#���}��B�8n�����S`;�^b,Z���,��%Q �x�z
�h�h	�v%Y�E5�4��x)�$�bޥf%�ô�c��C	� (<�Nm1.q]�%4+U�`5g���Y�c�(�yz���J�VI��q��5�¥B�;�UhaI�}�c���v����2�V1yd�x��8p�ߔNh���J�������~գ��yēw:8�
C~���;�Wߩ%'�"xm�m���!if5w����u9�$E��ㄆ`J.slJP��Y7�L%�+:�i`�g4T��c�F@ۋ��E{�7A�))���^�����0��߆���ѷT���6 ���������v��Ah<�?;��t�����l�	���p����\%�.B/�y/z�����	jȤ3� ���k{OQf����w5�sƶ����k݂d�7tF���:�M/)��a*����:��5���B�����=�@��@�6��A�)�wN씜ݥ~s��\���h�]�EaW�
\�k��T��Y���D��ܮ�F9#�������/��/��X!��_�ƛ����0f1��$VD�5�=�~�JƸ׽ٖ3��>'��ѐ�[���hR����YL�t�wS�0�L���)���+1������?D.���}���-lI��6�qݨb�2R�T�\�y�|�I�m����GxN���,-�~��(��� >��{��2�������i��C�!͑;���U�/��m�\��P1����)�H��o�, 
<)꾤"](��UIt�I?��2�jd_��F;����P���|���
��+l��<��0,�FvT��=RŃx�û�~�Wf��!9e�-���A�B�����ߛ0���0z�E�ԟ���q�@uX�_�s�5�g�J��T��{}`*�o���+80��b�(�
����?�%���T�_ӥ$q+{z%yy]G�e0�A��F
���y�D���+o���b>V`���X;=����*9#.���+�QǍO�`�sհ�IO�D��������vgvD`��ōe��G���h�����4`�qh��a�XV�n���Cw���en��fG��~TU@����F�����%�V-WUoR�,\�9h��e��,�����Uf��|����,�w��+��+�	�Qa�W�Y�P����T��JpK����Iq�6,�/}��ڌ��mGKM8�¼l�E7��K��t�^��'�Q���/�w��"7;V l���H��a����Ai@)�X�?"yM:���DаNX�o���WaPg ��N���.H�����m~+��9pV���`I`N�պ5�����p0�jW6}�������~��n����p�d��+b$N�j*�u#b��VIpB ���Ϊ�%�b?ce�0�K�m�״Kf��L��Vs�=h�������~l�z��0Ls)�ի�����c�]�v5����7;��A)�t��j38@wohF-Oy��B����Գ�;�PvnCj�����"���G$��k��=d3��H6C�X�����[iR���;/�oE1�\���OI%��� ��+�>I,">]ea�_�j�����3�+IX���[�.��]�$w��N*�5/�^*;d��дF�����LoϷ%�|,8�8
���ӎ
>F�l�w&�S)��=��|�u�b��b���W'v{���c~�O��
SA��R���Í��/�~T�B²��=�j+��F�"��Y���E�ŉ��^�8��q�^\*G�f��¸�㵻9vy�1��y[f�՗3��;�񝳟w�� �0��M Y��hD���2ms�]������Ȃ(׈7^�,fd��o�3}ݚ�ݾ�Z���9�cSq�iE���1?�s�W��]�f.��኶�D�y��g��w�������Q���������Y1��-�7�y+�BEn��^^a������Jީ��-Ey�=��̯ܺ�8chp�\��؉U���t�f�М�
Ɯ�ҥ[���Kb�?R�7&,�Q��^P��my�?(�* c=�2$E�B�s��LN
w4��� �v[���@�@1�����ղļ��:K�-��|�>˘0d����idO��od[�%��-�T:���>>U�b�R:,Qq#�`)Ӈvn3��V�A
Z�C�;;��8�?&�h���L�~uX�1y�G�Guєj)W�Ƙ�:m�a��������RX��m}��$�}4�._w.*{�- �����E])���o�=<��:��f·c�����\x
�f��)z�7&�J���S��yԅ���  K:8&c�Hl�t@��c�*���	/�mÿH���r�	��8W�<�-��>���n��+�y�{�n�ݎN����b9�i�;(4��#���fT?9��[���a��a�l:I��U����T�< ��Hi}��]W��mS�&Qsk�V�V�V�
%y?�(��G �r1�վ�&��i�JC(O��=0�\��>�j�e��/߇�򽣤b)Y$���̷E珥B,��&�~��gee�����'RQV�oŌ�Pj[��G�R,�;<��ǆ	 i��(�Ƨ#m̈.;}�J,c�!�x[t�ȏ����΂H(�Aw�uV`]%�p�����~>�}�u����D�5q��nI�� �mW���!.���X�5L�2����O._�C��Lɞ5�������k8*��w	֖�h46��p�|g1o��'k��M��ȥ��9��If�M��;j\"� fg����h��]� ����r��6Y��;V%�Y�1�^�C_��W��ʼ��
���pq=7�9j"��,�š���x��B���\�����R�Z�&h��@r�!�q��.^?[�lG�=��ͯ� ��>8ఊPo!�mţ�>>	u��,�����14+?
�C�
,u=� c�I77���nEnȰ��3�����1~��ש��C]f���4R%��k�v��}�Q�ҍ����S������@��'ڃ�j���H�'�
��`�2���0Z���b/����Z=:&7W%R���o;�+�)�lWxD)�ȱuY�'P���ځU̕fh�:G6�a,B&�KmE�R�����!))�kφ��>s��lDv%��߂��O��ϵ_~���|l�J]�]����t�K�k���'%�]_m��������\�s���o��ek���D�����a�T� ���\�!&G��/hl�Ԡ@m��Z4����_w���Odբ�zd�)�mi�C��r��Տ��LbQ��h��qφ[��I���8����\1-��v������M�e`i���ӑ�p����W��$�<`�"�b�E�t[��W`���}���m���%��������[�ٛ
q�Nc5'�{O�W�s-���ܟ6���=5�tGTb_��i-��{���ٚ�,��+�R7��Z�/?!V�KvCA����?5y��P��|�f#W���WNU�/��E��7��z��~����"��sf���T�v�ܨ��/~v����D#ֱX��&̒WA7�֪�hQ���8/Ri�g��[]�@oFN�q'�vzdj��_3ib���}_��m>��	)�a��r�R���4�kY,���u ��+G�zQ��D��&%��c�~�[��!����z@�N�5q��~�+	�Q����[y���fa�9U,��M䱈����_x��1�����{XQa���"X�?��5"�Z�.g�~�'g��y4�4��gǣ�Az���s��lA��{��������-rV��<�vd���q�@~��+Lǃ�)�/V��	5=�3��7i1!0ϻ�]�FQWP}WP��-C���G��.2��N��P�^���r-��KP�S�e�ڼ�U���Q�@b:a�K1ifʡ�Z֊�93�=�pZ�*a��?��Վz/Cy'�C�R]�b�(�y!:l�u��Q%y���Z�кjR���S'���^��6���=s:KXi�P�m�|ǥy'�G��nd➓���WD�&���^�^bb�Jv�k����߅�eH+�׻�ƭ�O�ا <E���v�t])��պ=��}��x��Y���h?<�+*ϢŨC�G��md��Q`m��I���_ ���4��H�n���7_Wїg�j8���`�=�� �}����l~�gi�yw�e���,����ʺ<sF�����u� �����n��k�s&��e�Ƚ�n\�[Q�Ó��f�O,��Ꮥ�w#��C��4'�G�vxU�d�}lL=
j	x��3YS�&v�Lo7�3
Q�F�8�?���s��Z4�O7A�}����8�چ�}c�!�q����qr�zC���x��m]�	Mj���t􀰽n�sCV�O��v�ȸ�ŗhR���M�>��,�<%��6��T�R��c����h�@�^�f�7F~�~#��gA K_*71���?X��e�F�#7��W����a]A��|k$GN�.�I<Z�R�cS|�5e!�¾�����M�{yH������F�L�����׃�7��~ ғ�_H�O�q���@�$�����n�KL\������m��&7�˓���ĥ����7���A�����mb��&�,�Ǹ-�9憉c��q��߆t����1 �����s�ۙ�m��iw�scq=6Q .]��t��ߚ�B��T���E+�9N�sv�Kʪ�U��{��������$���59ƫ}�s�W=����� ߻()axy�r^U�F��@��Oo X�@7�I���0��mZ���Zu]sā⹿��_oo?6�ɿ��;dj�o�	\��z����X�<&���ב<E_�9QQT��g�"cȼȰ�� ��u�/ (f�ݕ��/�@��ɺ����-���i��6f`̯��� Ot��Ds���`��+�ڰK�w����a�0:���CCG?��e��V��ć�qx��3S�(]�] �n2�a/�sΛ��)�����P�����.
���.h���v�h>Ӓ��!(kq{�ZC,�ҥJ+�F"W�|�pTL4p�J�x"b������k+���������^�8��2S�-����WA(��`����N���Q��K���S�h�a��Y��r����=|���M�@C�y�o�>	4�N��KQ�[�Q�� ��ޒ9��s�0S�u^�9�`u>�6�K6і��A|�A����jޑ�O(F����ʛ��@70��Q~��b�W��PEh�Ī� ��*�[@4�r��N��%��Ӹ�5	3l�'�[�`�K�N��J��E��4�x&D�*��7��(����+A��XƧ���(�r��v���|9���p%|��+F$_-P1�����,� @w#�gd�=�{?�zy�<�:�_N��x JǴ"-%[�r#�)�y����|i*��t)i�bәϱ���t�	��D�I��gɎ� ]�rt�;�1��cF���V)51����g�����8*�,z:����)n��Ip�i�']�X
���u����1�P�HtZ_"<�hh��?ּ��럋�?���M�Y�v�_�XE�_���/́ڻ3��b=lsdL;ܻцsI�D���'�χe�G�R诮_��Y�c�S��x1�g�������~I:��NJ.OG=�����^ľ�ΏHN�,B��I�l���r���V��В:���q#x��ے�ʊ�d3\�Z��նh�'��Q<pF��^��wR��>n\��p����űt׵+�C?�;�Q��1�]�R�#���w<:%Y���C˶S�K�]�Q�VW�#�3���)eƲ|GsH����C�E]0���x���=̦�Z,�m������>��W�rJ���S�ЖO�/F�����iqd�>DsQ>��T�t�����t������G�\+���.9(�t�ų��
��0�٭y��"�<�J�&-A[�g�L5P��|���@(��k��]����[�Ե�v�2	�f�-�8���5��s(,�d��������ܹ���cư �v�>���8�Z��1��4�����I�R���n�4a#�U~ׇ�w������ֽ��=�3��̍Fl�OTk�p'^f�O��
�<Q2�Fc^�P
�-�Jȼ��t�G?x���V�"������[j�=�-j'R���},�ձ��\�DcIBC��Y#w���9����ge�N+�Rj�6��ۨ�d���B�G�0�;bN엱�-E�eRƣW����� �"t�*S��v�w	�iJ>��l]�]�Z�ϳ۹�)���2j2K8r��U{��<�N�=s�Ճ�`�;�X�II�Z6+�ě_��ꤠr;+������.�Al��)�7�d<�;{ bL�zj!�2W��o��˥1'>��`�va���	���-�&
�5W���ܠ3�`���B���Gp��'���/^~M�aN��lwE��T�*Ot���M$�J��3]�0d�+��XY��QDDn�1�T`N!�����P3}�@������C.���h�+�g����ɏ�������+H��.��Q햰q"�7+�n
���z�����T���#�-q��F`UbakD£/���\��b��8<�I"y�R+�?���sq�+ ��z��Gs�����OΣyb�h��o����:3s8(��m|��kJ��eμ�=�0����ψ���� a�\��#��n�n��E��9Ŷ����p��&K�:|�3!��F�A�V���7H;��d�U#M1���}�OJ�ZA2UR�ݠ�v�v`��������I9^��[�I50�ZU^�5�,sS�ugs�_tw$Y�9��F����N(�p��Z�7����J�)]���3����	X�	�^�F�ڔ~H��M����T�<�K'y���X^m�SC���_��J�5�Nvyŭ�4��DK��ܴ!�5BCUM��rB���d��V���v 'z����[���5;',9��7!�/��-?����v�q^�-����Ͱ�:Z�-���O~�ؘ챆R��k�ϙ������__�f�W��u ���wK4���Q��y-Ļ���Εԁ>ΕOy(�4��"FK��-�f����Kq���z�f��E1s�1���K���/}�"�׭WԔ�K6rMtR�hZq?�	�?�D��;O*g�KQl�D|ۋ�wy3	^{!%ީ��j����8�_ڲ���j��x�Yed!�d"�f�{��e�*�L���]�f�D�%2�8����s��[X�J��O�V��l�$�a��П%���NFj��B� �m��1��o���~��*@����喈6m��vd���VX9ܠ�@?<�1L��u��?�3��\ ����t�a�-�j�H�1��a�}.�#�}�z�Ia*�lYP1Z
,y�q&�Z���G��{��@M�w�m�@�r�J�o:�Nâ)��VZ��9#N�4F+���s�$�6��.��W�ց��${|����}В�PcUxnG��~�U�/�? $r)@�#'B�� vWPB�1#�Q��}�Gg��K�!�꿃&��y��"��@W/�1zݛJ�!�ޓ&�F�bB��^�`��t͎c���nL�l��~��e�g��)�V�=�G���n0�4��C���O[��/��B>�K�oB3���k�A��qi'�ʑ�����^-v��[���?���j��c�g�༌�[fz� ��N{�62Z�;ӕ�����!dUJЁ`��d+�Eg�o-���M���ی��������&|>�;��P@�����M5��)��c��4j�����F��u(ȕ���\�\YG��d������d\�1��7jײ�L��ӕ�m'�W�I��a|xAl�� �ZH��R�:�My�Ӆ�Έ9�w�(F�$uZ��=�XKf��K�B	�c�n�d�Ϝŀ}��Dn-V�av�ep}����z�W�-#T�-���#1�y��)&
Q3d���Y�5JE�(7��S&�w�q(v�U}�(����A�Ns��cb������4 �v�vɊux��X�޲����6�G���_�������s1@��w�����t��^*���1`Uy0�5z�XRA��b昘yL��>2�ݦ���U��n� .�;�
p�8zYk?PM��{q+Hx�P�S�7�]*�˥�������G]�s���cS�?!�p�̒=g���A���kC��k��vMH�����%���\,+iw�h���Y{�-D��V�c`���rwv�t��R���;G3�d'�N�{8�l6!����Z��f9���1Q��#��g�,Mp�]�	W���K&�1�'Fas7ʵ�^���'��;^���a�s�oש{m���@���'�w��<n�d��)��݇G]�`���m�5��S�yz��Ŏ��!}�JO!E@AfzY�av��8�&��툉 �}�W��#.�6V����Xٜ"IH���,6��/d��  i+��́k�+����>\��2�AJQ�|&�Y��^��M����(3���e��K���7��bӝN�~�cQ25�h*Y�?�tʰ�n����MT_@��k����{�,��Կ����1s�V���H5U���8��#�99�������D�C��#��Lɷ��������\Z�Kv���ʚzD��u%���|.
o���<����5��Q�����X�e?��)f����&�`������7qR��l�J��yW7��*���^q���1�?b'82����P/���o�>�cDʾ�����ֻ�6X�/��(�o����.D���o�9����8��0��n�3R�(޺sߨ=�.C☮��k�z�Cn������d����5d*:a�2w�A�hr$mS�����nQ_ʾ�ucz����p�]s�VH�V)��w�Z���^9���JT��B��Z�y�J��W���5������G�et�i70�ng�[fpm�����;���sQ�$P_vWhn��q�S`߱���C80��ͱ��C7�%i���Z�?je(�*/��e�l�P3��)��aEM�6��;�B�!�G_��fF���F3e��C�tc�a"���=�ݾ��g���{
�+9+�.Y,������/�j�t�,���a]�ڏ	x[}�B���ZC	VT�d�n�P«�ؕ>�>�shhh�܏�+��ee�]�9��]^���g�q��k��,oT��?����ft���m,��W
뛍V���3*��}�Z	 ÿ�=��)��》�9lQU��&�1�]z�?J�/��h!%�_�%�[������~�����C��<����k�V6s@�-Ѱ��N�+�Ml���01���~1��sF�JN��3�H�O��(����#(����"øS����B{ �*g�@�L���C�P>���YGd�t���گnSqG�&���J^6U�_{{��%mP��f��^�\�pU��*�Ie5V����K\~e���p��w�d�Zִe�GT1-��ɓ�svx�պ���l��Ο5q��]�%G	�&Tդ�Q���w��DR�:hKW��ko߻�o��SPg|j2�#8|���#V`��Y�ڈ�!�,u+�@�=7�ܤ�C�>�*��w�)�>fgد4���$�����;��/^��ѳ�V��?a%T.��۽�B>ݪEI�DQ�#��f��\
�: �V�Y%W6���4]x�>Q ��<�jIB*���)mP��F��`{y�X0u��Ш^����j�c���,� d(�xd"#�\�w�Mϥ�
"ِGz�ۮ�f�%qU�S�,�v���v�u�Oj��ܻ��=A��٧"��a���� ��MW������ń��u�c��%P��E���O2Dca�
J�M��*���ѡ`)������J9ȕkc��S(M%3w�K�d�A������^�ܿ{&1�K>"�
��9��?%�ky�ۛ�Vʠ�� /�9�*0{V(z��ᣃ#,��|v|xss���\U��DeV��6,��D�!i7�l��b����`׌��\o����UwA�θ W]z��}`v=��6�h��&�s�߽�=E\���̹2��B�	�.����dE�
S��6��G��X���s��6a�o.�s3�F<�a`ˡ�^����|�ė��1G���-�F�h��\{'M�3�+�#�U��'����\�5�̫���8H0��Ct�.��[�J,r�L�>�T������C���HeD�<��6����b�&�.���k���ZB�Tiw��e��\�T�G=�r~�����"����n&` ,`3�Bj�����i"�u����	f��\�bsb�N�k}ժU�􋆳�(��e8wh&j&w�]�4Z�kxv�����	Of�������0^L�_ğ�~!C���h�!���z�6��өd�NF���]��33�!��_2��l�y59$YϪ��#%jr������� C�v����yf�24vs��R�~�wO�ɱ�s�,��'��t������-�����9�ضb�k�g X.��p���6�k�1\�z%����zx���t��-�z��%5�8|�M7 �C%ze#2f�`��ʺ��Xt�(��@ ���Sb�F.�;�[�$�)n��koW��{���<11����!n�;�t������ ��(n�����$��}��+;�	+¢���{8�+��2 qR�ZX| �Y��p+���M�|���y��Ζ�eb�,r��B� ��x�N�O�d�ns��g(���y��׹�Q��f�����/��f��	��6f"'y%�b����J.��t ��B!Y���\k�2t�Ӟ$?�>�:��f'C�.0�t�X��Ӧ���]�_�r������U'�K���;n�h�%U�G��-���zG8�8�i���0�$a�8ց�&��%^-}���q�*t�0�V�y4M�D}t� ]c�9�4��]��,G�ɋ����Q��	��c�8�ԅ)c�w�{d��C"�c���M�l�����	�M��|i�2�#�fҸ��r#7�7j↸e��W�f���5�w�4
=�8�����.R@j���̡E�	��J����oqF�<��4����}.2�P�t;Lf2�7͋��=�#��Z��נ�1
��,L�o���胋�:q:���?�k�SCS]�DN?�&��?g�˿E�p�r������#g Zޥ�J*�p%}���ӏr� �6e	\��%U{Pr��HF$Ri[�?�^�]��1��J�2�<�xu𒈒��7c��PcJ�&��H�߶��+�oy�>1�&��K0*87���z
��2��҂��f_�ty�_7�oQ�]�r� ��6'�LE+�<y���)��i(V�>k��6Ԧ�~����LX@�eB�3��#�@��9e e�����,SO(@G~�"R��T�"Vk)�\�{1��c���;&F
�ß��Q����f���S=�]�-0�&l�2�;�HW�]t�r����ҋ�pP�'ҳ; gu��Z؃ˀ�cQ���6�z�H�����ձw�����5�����^دN�|��.�я��&�Sd��L"cd!^����J�����Ty,W�q͡����4���/��T�yՓ2�2tjd:Z�S��|7Н�P��ӗ��*��6�%j]�r{�t$y)y
7�;��Q�1���薆 �
� ����v�M�r@Ֆ���&d��u��}�q�fp�G�6k����eA�FVM>�`����I�}Y�;g%)�qe�DCd�Sg�0Jc4v��A��0VP!||�}&f�¥}�j]�j��uΡwI%]�����)ET60S�T�J��i_��	}����C�J����i�"W&HH"��}K��,�����-wV�9Q����{ ]}�]:���#�TdZ��1��m� Ns�Dz��ZښKZA�*�RUb	��P�$� �1��� �h[
��'�M[4�������a�f����9����`ly�!]���s�,��khA�2XâYk2�I��°'�Z7H��ʞ5�z	 o����nn�%.��^wGXƀ��gz )�b~ p},�{��
ky��0J� ����x�Q��)�[<��$)NX��z�
���|
_��vs�y�ET�1��K�$���1����]�)+o� �[��mm������nr ߽8�ShL�=��@��S��zq�Z����jwWBd�X'`_S�׸�9���Š���"�g�'����>���kl�{K���t�f����T��K�<~�)Ѻ=]��
Q�b�B����B�f�}բ�A�̭�`���s�)��Z���!�Z��!޽�l/d��� ozg�J;�.�1��2�;~4�s�^=�����х3hy�q���>���1�X�\�Co�G_�u/�R ��j�O8��b�,"!�c�j&��0h(�YRk̤G,0�k�����	�w���_e�8�}�lUI�[����OI�LOl���K�%��0�^���p�oK�O$���hs�����r�7��=��_�$�����-ƪ�C�6��fXiﲋ�?%�Y�x0�H�Y��0{4�ڭ���h� 鴙ѐ��e�uB��A�T+ƩYI 7֜Q�E����>��]�̛d��9�B#��s����#��x�F�gY����<c�؛�S���N�+,m:�;�YN�+<��~��-嘪9�X<Ed�t��$�Ap��AR���Ѹ{\�:��N��x��ri��PHNG�~���"���Gϻ' ́9u��ok��&�f2?��x�r�d:�Fo}q����?CM�"���(��Z�8��N��~���Pi�X힋.��خ�>7�F��B��@�0na��Ɋw�� 1k�YrZ��`�X���̍6LW/N{?��Ag@��}	-���Mņ�ZjØ3�I���4y�ZW��J������Nr	�G+��Ӓ:�#����tgl���ݤ�u�$l2���Qg��{�����ᛢ��
"u�"$��6w`(�|| ������*ˇd9�- ɐO�4s�,{( ��.�̏C�$��0��~O��*Q�s��
ˆE���+�
���`���/5�<i���>��#���Z�@i����)!�r���ˁ��!��	�V��1y��m�b�B�iܳL�Un���u$��nK��Up>�����x���QO�m�M�d����*%(�{���ºl;/�4��eb=����!ޞj���UB�r�@w�u��C���;����۠�WmZC9���@7���D���'wo4���G+���g\3�;��؈�B+�:l@���VZ����a�.�y��~�P�C�?+Jc�+��8v��U(�˘>��&@��%*&�`w��K}�4�R��rq����)3:�� �.?���"�7���5S��
�� � v<`��M�N�\��P#`�d����������'��/۸[vϯB��<RI�� ��2��	QA}�Y$c�>qY��gM�~�#l<z��^e��}���u�Aax�-�$n٭����y�\��I�}w��'7�����j�k
���x�o��<��+h�K��/������K����[8���=j��p/��4��X �
'�gRt
?M�;
��jY����j��&��)B1�o�Y��|��	?UM���aAK���A����l@	
��������wH�_�DuG	 ���8.~\UBm�wyC���Ĩ�g�b�y�Y�o��4[�cr2|Q�"��k�$�]G�&zB�itcCK����jG-�#�;�j�dL��M.K9�8S�����z�q������'�L�,w�
5�ؠ�G��c��Z�/��\;WJ��8Th)@�o�D��%�H
�ƭZ�s 8AF^��$�Xy��?�rT�q���d�5kP�!=�%����Lв�4�P$�����!H�7ɘ��J�D:Qzhi�o{�&�a��7�Qp�I#�N�W���:[~x��m��[��s����F~����g\+����Œ��&i��z�G�{�"k	/]��`׮�5l�gNܰ1�c�Y�s^�8�}WtQ mNGP�N���f���;;��2�D�k��K(
��W?(a�^$�7d�P�*�|��z�'8b����V/]4�UDe&ߚ5�d'GC�#�g���z5�-��T��'v,��C\��� �i�����d��*��m�d]�)����Sˆ9������2J[*��G�vrp�4��za�`�c<��ph)��7\
����s�EA; 3G��O����2[qE7����g�yGo�|u4���]zع�����>�#R����!��=P�ڌ%q,�s�t
}3���=��aSH%�k)̅��<"D��^��a���;͆M:�uLs/A�hw��%��M��H/���_לt��h�U�����R��Bt���}�F��K�TK��Ɠ��(H~|��1L�ϝL���\A?^����������]���1���)�x=�1}�:52���$�����R1�K�۞�$�=k�6�qT瞩&��؅ΆtM �\ķ���Q��L���&~�w�g�9�v�tj;5Xµ/X0c�ֻ1�371�����՞�E��x�6�~��4������E!7RH]�v�2��O�S+����(��2W�t	��=�0���h{+����[�F��jk\ H�n��FJ��=�/�Ds� ���y�{��k)������"^�R�r4{.��,{5�Vd��C�@Ŭ��L��	0��(�a}����ا�Nk�Lz	!��X.��l�ݱ�ekRQz���*�Uø�A�尟A��BfC��͕,zϕ *��n;���\_���E����z��?}F�{�b�^��F��z�"��?b�q؈-Fr5���19M�L�-*
������+���AL�<hmr�KS`�3^��5�RCa���V��k���q�����%+!�	�|3W�|Z�đA"��\�������(-F[��a��Dw�Lo=�[�����a�����xfP�}W��]�(9fn&䂋�J�~㛛l���+��/���*F�|�^L�O��"�������j1��DmH�����C"'��8��:��Ր[!��o�)z���*��A:�Ң!ޜQ���7���S���u����r� A&s�yB�D�^�D�9{h��9=�?�1��5oe�:�m�^�<��@���)�rB�ғ1�v����#�V��N���/,�\q��>i����_���ПT�rk�|1�І��$1N'F4w{&�:/^��M�ߺLօY�j��mh�*�ϵ�������<q�5%c"y��+bީ�fm�3��/�w������zw���Ơ�ԯ-<Y��+��/(�����U��3s���p�m�Z��[q}c�;x���'��w�8C���������C*��l
Gq"u`
�綮��a�}��9	�S4�Ԥ�m�1����蝋FT�{i����p�9U��{��ƣ�I�7�2���I^��g9�P������щ*���˧nx������S,J(wTԋ�����LsE����Xк��
U�½�)�xfl���J`��2�F�:����X_�X䗕:Iqj_�{l�Yѹ Ծ��{ѕ]��{��!@�?Q�v�n�Dg0K���" ��\�C�ն�	Ua����'��<~��+�����cV����y\���¦U�g�7פ�Z�-���}�)�ч�"
@�J�n�L%6�����W(1�+j�1=C���C
#��0�k^�W�����?ŗA��9iT�H�>o��ق�<��v�
w�6���M���l����"�2T�Z�-����)�^Ls�QSl�R�$����G����7;��[cA�0^r����@[Z�^s/�$53[7�=؊s��x��%�2�/s�����CY�y�B�|��������S?~����g�q7����,�]�}wH����\�Oa��䜑��ɫb˹�d��h�R�Kv6�E^�~p�e��n��mr/�����B4b����G�_�>@��lⴻ��	d��Ji��!6x������Pb��ީ�\�B�R����I`o�ѵ��]�o�m��4�8�0�r���3P"�*��ȏh�4J���+�M/!���V3�4�+ob�
��q_�H6	0���������R�8TR�S�P5J� �ZVQV����#}�']7���ɷ���Q7;���3݂.^JW��Y�"b#��Ϫ�~<�bE�����$H��m��r�]�*�<��q�q��E��BLC�K���{��[^�������c]El5NJ���gx����X�4YkS��>���'����
r�`��[V���5��rk�!O�ׇ�	K`Nj�II'�u��$"���\DJ2B�5i�lư���*5���܈� �T-�F�{�жt\����F�~/��m}��;i!������NHY�"�����,���;J�\yU[B���ⒶR"V�k���C�u��IҞ���!%�OD\��|���9�#��s���9ҽ<��̗��t/��rk����b�mh_��A�-�;��UG����e�~�������۰�oq���邶뚏)�����K�؆Ff���b�<�Ќv+�]V�a�L��{��|���HՓ�yd9��a(7t{PIJ>j�s���{�)bO��[bJzB±Z�7{�	���QG�$7	��	���a��f��h:�DEe�����������"��)8����C:n�U?�;S8��K���O��!�M��%¤��X�݇&��'U�d�8QW��G������\M`��*ؿ�ڃ�!��܂c ��3��a��D�v�m�)�q�a6��s���bа����rgJ�/f�2��@-0����Wq�Ca����d�RFI^1����p��'<b�����:4Y(˗-����\G�&9��)qҮ
n@��yMD�k�s���nK�I>߻Ûg���`�/FVP�4/�Դy�)�z��$˘�(VhG��d��9p��uS�EnKD���1����6��P���/��^2͋���"���S�I�_}�I��HU!Mc?c�x��� � Ͷ�AJ�*�V.��W:O�$�ʭ�����z�Ծ�>�CkB77M��Epk�:��D���-�_�dS�QKMy�;m��T�Rp���|tLv���>�̾<Ug#� b���Z�Or�ۙӢ)a_�˃�Ɣ���o��R���E�ن��v׺$�K��uE��?4����^n��I���/h$p ����z={�`y�*�SR�����K��م)��]�/aw����������i�~���B�jυ��)�K�5�b`�.9���n�/���(X��giX���UN<�#�Iw�\zӾ�v������t��L��(�I��ԱҚ��:��p�;���1qiN�VEPR��w{���E�ҧ�Ĉ�(�<���a��qq��B�d�)�t��'�bX�2�k��
�Χ:�w��0k�1lT�)YGE�v�s�l�v�Vn�����WX��J餡\��Pܣ-pS}���7U,>�<�A�r;�n0��	ë����Xú,?�=�}�� &��W��;W}}j���Z�Ȇ�C~�^��v���<��g6U��h�;��>4�L�����Pɏ�1.B��<���AQ)��z���yZ5��>�o�A{5��^R5�����R�O}�/��m_�k�_���Q#�E�1�,��:��՝�[�,����?A�1���0FT�֔�`��>f�|���H�%]���Hp-�T�Z<�����YZa�4Oƿ�νR�)���6��)��W��
ȻH(�_@�*���c�qhC��[is�rI^��q�{���`�6�ޛ��꘍�-ܞ���:���Ŏ����#�>���'�������vՌ��)e��n�l����+G
+�=��k��!-�a��T�V�uM��_�˫���΋�\�2a�|J[���\�Z����39�6�|��O�[�N{G��?"�	ɪ�qzȺ�M�eXD�'=�cJ�]�����2!zu"�K�㚔�1P�ZQ�Q���s<��01|��(��бH��1�Z�v���!N"��:��P��n�
(<�3r��Rw�-����۝�*���<��}2Q���OĔ9N͞C��$�Y������h��9<��)�nA�by��≳�3BX+�Y/[�Q���b�E��:<�z�E�Bݒ��cI��#=���
�+�Q�&T�o'ifr�8��4.�KyG�^����;���ٿG��L��Zk7RG��3��������;���]lm���4wTm��ruˣRL[C��)�����<5m��(]$�M,F&�Y#8k9�r���#l�0�#}�� -g�,�g�K�t�I.���Y-�[�<���X������� �
�a������C�n[&bT��jao0B�J���oII^����	&��X����j�W!���$����8U���p����v[����o~�B������*cS�A3w ㅂ��8�ۘ�Ô��+��ɦ*ҸMO�H�}�'#}�0�jS3��.Y���Z���hH���!�滨�2,:#�@ߟJ�O��x^`�i8�'�&b����!�
���T��\�V�$ �DVj8|6�D7�F�8�~'�L�x�Ts��|'Ȉ�ۡ��;b	2 aX5WPv.K'���V��9 ~����;`ߛ�hɏ����?1��z����C�׾r���
[Y����R4;ȃ���0��d1'��1�wD3���I��T���e(�$��r[%y�H��8
v_����T��z�"şJ}h	�b[��>�ͬ"f �!��@v�B�����e��C��SY½ �2y�qݶN^�$�)��咺�q�ǯj�<m�/f����*������= 
�{�ˌ�i\4�q[yL5�H���^�ٓ2s:YR�:U]׫��Ͽ��v?���0�t�إ6E�0���zp
A�Ɨtc�~�RS�t�[��(��T�0�1��l����ҏ�<�~�r8#�-��7V	��?x��z�� ���S�˺��y�����"<y*�Ø�\p6u�eܥ�������r���I�G�Bѽ��7@��6�i��?y)Q��P-��u���g'~�����
' &�#�Q�4o�� }��ҳ�^���MCD���;������/�w�R\&���Ma�6�T�ĐS~b�V�p��A9�'�W��!��������8����r@����	6�����_������61�T�E�kFH)"��b��KnF~�r�� �~r)NN��p��{J8��XƓ�s�N� ҵ
����9�S]��;x7�zQv*M���2r���ȹT��zB�μ��l�880EG.p�xn<5���?~^餚��ߒ8��X��<���B���i�l��'6r}��q��\�S7A޼'9�i�m��oD_����J�&����y䮜�z��0#����?����+�Z�>����m�Y�]Km�`)��:��9��)I0e���a�n�?���U���.��c��`��_i߮�� �s�%G����*[����6���-�Ɋ�SמI �񍴰gsz�^���I^�����P⢐ӌ�(z �	��us:�.�ڴ�'��N�
A��G��x؏�d�mh~O&�pQ�:0�;8�#��E�"��4�D:V�Q�k΢0�t!�Fg:��+�5���BTa�t�]]@# �R��{DV!��t�~��:�a����G�u�c_�q��f��1�ή&����0�B��ā}c�y�H����R�.quZ7G��b-W+�3b��V�ֆH@�����t	!H�2V��LXY�7��K���[5��Zf%j
^v\U�5	�y�>;N�,h��҈���|��o�Ɣ�1��4}z��&Y	o���y"���Ɠ��������F
�܉,�4'Aָ1���$۞~}НңǍ�wLᣳG D)]&g��lf"��~{��-:��|\�@����n����P����Y4�i'eA<���OD�O���@�ӦNع��5x
>%�������.wUG
�)�{�!���0$�r�0����w��T�_�sse�<����t��#v7-H� �xAuN���0��g[5������(��5G���].�7%F����_%v
�~S��1�;.C�NG*\�ӇJ�m]���K+{X_�n�l�WD���{t�ǘ������nQC:�璶}W�a	�-v��Z2C�����f&ha�	�x��}g���q��0���"���eq��t
���G�vb��B�b>��.��9��@!��@+!� �e~���\��%k��޹tz{�a�^��? ��h�V��}Jͦ�t�:''!a;�|�E��� )���ӹ�WA��t$IT��"�< �vU��a�t�2F/֦P���Nn9;H�#�&l��_:5]f$'!�^K���F�VA��E8�N���{�* �4�!B�� ?h��>�D���G��[�xh^vġ�;�SW��?�H�5�����KYK枹g����A�M�[��� �R(��5�2L�{��*Y۔D���Zv]����L����-rI�wZ�*�ܵ1�I��~	��'�O[S��@�9�4�G�7p*Z�0td粌�锂_��g�3��2��g7bK�)���ni-���OaJ���E�[N��yӺ@� ]��D@�Mѷ.*��u��a���}��[BE���v}�s�KB40M�!�V=E�W��Ǒ.��.��ڠ��Ef�wdr|�B��R_���2�����m��h�c�%�Z?�߉���
�'��u?�y_S��Inڨ jH��LVn!3�B�pX#�M��gRx���x��s�~�^o6�h9,=�����Z'~��,; �b�|+�ǜpBӰR_���I�a't#��)��4u���1S��.��~4W}lY��L�u��yp��RT:ۗO������@$	0Ln1|��au=��0Cm��d��L��c��lE�Mp�f�x}�����Y�Rz�m6��Tl�FLM�T�v��Vz��*�ib����*�W�0=SԹ��iqkQ�gbdվ��18�b�4�%�����aCЗ,%����aL�b�yVm�$vɜ���E<�X[1���s?���^�i�ɸcP���/�_���̩&����窏��HO(0�:�����8��Ŏ��bS���1�v%�؉2�U�x�k����W���mP�s�NIK��+�&3C7�	r��u�h}ȸ�SjH�N��WY�I�TEks<9���yݒy��%0�}r)�@��L��-���B�i�k!>k�,�^��	���]�����	�U���v���\�s�Z�'�%r�P���Ӣ�<���A��<���^&;��L�f*r��gɍk�oX8������eʖ@U���L_]ڐq:���-w9���Cp_�0����΢�Z]�Ͻ�!l�������������@�����w�����Ժ��v$\9���[G+�$B6�n��@��_��ȵ�eoy�kbe�yNE�.�8X��\��9 gn��{ʛ����S8��W��&k<,%�_��g2ޯ� ��>�h��Ǯ+?(	���G�fN�gיq_���W�g��4�Hs���b�?��ڰ�;
��('�%�����tw+�-�WJrk�&傮s,��s׺����sX��bk+Uz�-���������q���.�Ax۶�}B�7�{A5����Sڗ^��"�f!�C�J�f�+T�T�O��t��s3��q�T~�-�
.	B�7[���1��,�=�8P�1�\>8^�Q�he��W]�'���5!XG�H�+�掫c�Au�e�\�ɾl��� �k�'l�^*m���ŀ��"ʲ�R�$2o�G��+�N@ÝM ���x�Y�	:#�����t ���+�pfz�g �;yY���eU��&��ݽ����D�	.��^*���j{�Z	��3��z���Vv\~�{�1���>��."YZ�-'86I���lM��f���=� 5�5��n�b��3�dF��ƥeQ�(��Iҙh�������K��	����75%�B��J�'+��_;�������M4r������G���5���[�X��^.�;�k�JS��.��43���id�)Ԕk���+c@6G�<�ګ�YHx���5�.�ޙm��E����.���=�8G���ڤ�ȸ���q����Gf�R�Ў4�r�(,��mvtA�P�q���6{pQ"�i��)��؊�/�+�ɵ��-��j�#�7���0�s�U�C����7�q�|��Ŕ�Gb�B?&��
�!��,������{��\3@��:�SV�\�K���j������U�S���j��;�S���q�������{s� �AJ�>�lJ�r��=��b@F6N�ު�b�G�Ų �p=a)��M_�8��]R����W��a)�)}¦@�f��#Sv8��=�ӆ?救$_��o�U�$��W��q��t��x#�Ɔ`
�{iA�w���;S��e���uo�S�R�o.�1|����yv�2d��s�$�"�g�ו��c����. ��	LN�Tr#6j%&�TϙN�Cظȓ�*
Z@����@�U��i��E�X�b+����=�W�L3���;�.��~��zM��T��B�ێå��DW�M�iߋ+�������)�h��2hL�hk�q]@�ǚ��<l�m�lZ�Q7,�̼mԮ/�8(���j ALt4pa�b�a0Z�pAl��I�!�J���y�t�sy�hz<�P��Hyr��[����W4ZN�\�Jb�G���/U������0�|�~Ƈ�9�A+��֏#xJ�<,D/?�.t��}�?v�sM�n�����_d̈́Y�,fcx-�R3��P���-C�䘗
�����HY4yj��󿖝���[�%��τ/I�Tg%H�wS>���3�P@���a-�9���-��섴N��Ռ�R#�_	\�;�o'�B_౟��, �?-*�����N���%�8����F�qyu��J���h����Ŗ��BP���i�/u�$�{���s�%#���粳֠3��V+����flJ����I/Tϑjlt����3��lG�J��U�ĝ'�%�K'�P� ��(-���y��o�x�x�ţeˍ�阂3ji�01JPC�ֳ��%1^���oKA�}>ƅ$=�*6k���t�WH�St����9<ܕ
9��F_6S�O�q�b��\XO��EJ㈌E���5�mj�;���ճl�����yRЮ~���a����H�|K�$O������75]�5���Z ��xi��4*VTb[c��1��ͳ���I`���+*u�Zzd#�H|��^�E3y&��~����x��l��Vhe�'��N�Ui+E�b������>�L^֢� ~?=�kشU�R�f�5��F&7�����m;{g�͋1�U�	�d|���qez&�ɢ�&4�v��ge鉝�'��=�^�+�j��D��h5�OŤG���u ��:�l��}
ky�Ĕ���6�d�����s��[�W%c �Z�?��)-liu7��x�v�_����jKCP���<��pBHA����oh�I�ӓN��m�n���k�#���O�缌��&oa�N��ǵy�(&$ݝ��Qrѥ��R=&�Xm8k�SI*��K�-�����5���vj�J�w��w�
ȭ��4�u��U� �W<�2��RF}:��3?7N >b�_��� �2���K�賻g|C�E��K �w�����#�?>Qr1�y4z�Rf�����_7FP�9�T�@b�(U֛������zZ��L����J���E�W������h��^(P�C":�����9���<=p�L��!Q��fZ>�T������h�7%Kr�L?g��l��+��h�s���ML?�L���N襵T[����QZ��w*O|ҥ�-�X�pg����0d)����v"J�$y�҂���p~�u5�8A���H�Ѐ����C�q/��fOY�TL.�,
�:�_&��:��#�)�_��&�ʓ�u�,4�aS6��<�䐱��y[�X���PN�I�����O'�6P��|# �����
;����J�z���1�[�r$`�k!z�8�An�J����xy�&��Tr�y���m����'��y�Pt	}W2CSk!G�]y~D�V�'��{�R\�e`�=*�X���
�,)��l����J����Q�]��C���G�VB܏�a@҈��/�LS�._l�)���^��GN�$�A�)���X;�t�� �L��er��d�g
��x�Su���l����c���������
�%�le� c��6rR�`�j����>�~�����֡�K 0�Y�\aj�O�L�qd;�țĽq����+`��-�b{�{��V�A�qJ�Va%�&U�ӬB(<���qB{o��\o&J�hE�G��jn�_�X�v�%�.ӌ� ;<��v��D��;M>GH�ڔ�_eP_�5wdb�e/����4�%�?�_m������+�"y镶���iwr{2#(���c�F����IG�2|fT#�lb��� �0��>�9�������xZ@�MJ�L� J������IE`y
�4*�����$S؊�|^�7esh����@혇Zi�^AΎ�JObܤj��:DcSl�y�R�|H�󓝀}�7j�~o���yB���+�'�P��}��|�/�_2I�= �d�bg����7)��#����iĕN�Y��CKl�@{«�G����3��5��{w���쩐�Xdsň�n�5�@S�V���:�n�Դ@I�3-ہz䫈v��L�
B��{�Zj�_�ۇ��.8��j+��gK.��K��:���?s��_�D�6_ƛ����߲��|����č^�5(��p8���k�%$P�*��6 h'���X`���A%���ƀ	��ؼN�0�t1&�����֥�;_�2��?s�CI�0���p��vAXԸ�2�Q{���nv��0@Gv�U���ɍ��-�¯�r�Qa�D��0�}�Z�nl|�ȣk���rE�WC"MM�Y|SRrm�T�
N�-��(�Ǜ0"d^OV�$�BZ��E��PxA�y���R}�톴�2EB|x%� ���ip���Av����AyO��+��NRʊ{�T�GBGz_��a���6���������#@�\C�D��`.���������O��̱��mLߗV}����M+��&t�;#��{l�5؝{�-9n� �?d��p��9y�jDk�YaR 7)���&:��ƃP�6�����"L9i�]�,2���q޼�6�&��B�Q���?�U��T���Cu�Lè
�g >հN^S�@�%h�4�A�7�<oo׾�
������֖L���CMPC5xOz�<||����j�l�B&h�L�m�`��!Q�^;�"#��"���%.�O�|�����ì�D��-���*��g�A��.���h�]n%���@���{��5���y���X�O�ԯk���z�`�rqĜN��j��/F��'0G� v�Y�gn���_,�k��C�'Չ�!9L	zH�N��z7 �S�Jv�g��|���t�2;�g_���M��Be��� Q�V���2�$nߺbZ����,I6�W�Fp��ABɔ��:dN��?
Hj������IHW�514��BJ�,f����o��t<l�n������q��%�|��sQ��Y
A��T���AHF\}�N�S����ql��̚��v�i�@"^9\S��,)4���r����%����,���pn�A*y2�X��3�	3N%��;V��چ���VTt"���7˂~R��1��Ѣ�q�S�U�*:@�`�me���q �g�U+��d}ʠjh"��A�v���!B1�,]�W�7���nj-���N�����s0%��q(h.�~�iWG�j�NR�w|w w7�C��"LVr�A �6��rx�7����£x�x[���ÿ�a�.\&X�f堑P�m��2df���~�A�&f���70�}��G�>:%7E��o�nbkc��dR�����ӯ��Y�A�a���1�����7%���J�1�'Ze��k�л�������	�W�q�ez>�K�x���Ȉ�J�p�d��S�)��kc��1��@�!�_�ͳc3���S�n7�>�*Ï�l�f��r�>h�Õ��\�W�o}ݱ�r9�{r-N{L��&�9M j�-R����A���E�r���<|�*6�L\��A�}�Ģ�l�.��V�Z�|Ѹ�k�>v�_b����/�p`cY_#,�H��N�q�� ʠ��Q����.�h�;��������df:EC��4�}�ՙ�$���4�4���/s�^+r��T������?��
_a���6,n#��� 1u������Tk��ؓy�Mq�hp�R*;�ɫ�]����,�y�!� ����x��y���K��wtE`Ei�O�q���N�B|	)�b��xi�Ւ.� 5[hiG^uFC���Fޜ5���sv�+�S{�p��٢�Aͤ�!N��Xn��$��Ʉƺ��׍����m��d�D�:ԩ�eyz~\�;K����W�\Ŭ�W�G{�6/r=Y��_t��V��T$�oP�0^H�4�"	��Nc{���߶������sl �gD.�i��R����IDM�,r|�����+��!�8�v�oa��T��ހ��䨳bӽ�W�/c[ȧ���E�hE�N���k�M c�����{��T�3a���>Rz�)jϙ�HЌ���s�F�N'w�q���	��g�{qnS����F�����M}M����np���"Egީ=[��3�h�g��W�;����u�®zťw�.��|0�������
ύ��&0}jcVo��_�i���Ae�ol��[O�{��1g��5����ǡ'�{� ��/>n��N%ׅ��1_+�W#7Zv]a�-�Tm��/1w1�J�����:E1\�W�Ƕ�(dH�&q���T~º�4%�X� 9ȋ������ׂ�w/	�oLU�I
�$ȏ�Pl](F-�@Q:�9�6�?�S���)��H����Ǯ1K��=��H{�&N��#"�c�aK����Dq�$����@��Q.s���e��|�뇺�i�N~MwH_ϤqD��L��� v�^ޭ|�-�<G�����r����;�EX��E� �Pϔ�!�
�8;`d֕��#����ut�(��=(�T�dM;��Z��r���ُ��U���%#x����<��������x�&�Mc�z�hЇ���������+Xѓo�-�2=|�;}&+���Oݨ���!3��J��<�3-se�t��bLu��r�m-h2��h2�ZCXy
w)q��as�	C�+�)o*ʭ�w{]�C�<ɶ��yQ/)0в�ɪ�����d�C��!���|<9
�2�#,��H���8*��^Ht�X~�k����en��G��_�
Z����K{]}%������ț��'����{�vW�Pi�������c�N>QY� �F!Ǉ��D�k^XTuGR!D���hS`$�پ�W;���vT$l)wl�H�����K@����[��y�f��t�U��甠}�;�Q�葺{�3�⦯�8!B��������P�N0!�AO�Ŏ7�_O���#�Ut��5��\��0O��T8���S�qs]�w�+�ء�쿑�D��4ޱ�cp�/�?�N����ĳ\ֿD.+��8�G4��|�hu �/�>��H}	yCF�_�s,Z&�6Kt�ݣ^��J/9�=Ov���J��@�$}]�1m	�b@ʚ��5]�?p�p >��z'��ǝ*|�q*y3d,�߅lo�]f�9�Z469���/�Ո� ���n�s>��Va�2��>��DO��&Ϝ'c1~pN�~�wb|s�>xAT�N���bE��}|�W����F�y)���C~8n��k5A�/8�d���`��d�ޙX�FC�R��b"-)�U#V"M��
�G�+r�J�U�i&b�R���F^�<l�s���2�(��W��3�����T�b=W�N0t�Th��P6X6d���cb�P+N�p#��cn�6?8�&����H�'DP�Ii���ڨ�<���3b�mg�ty��kn�B�Q0��"{8�9�m.��Iu�/����� -�E�'-��٥�� �a���m6��9 ��_���91d]o�߉R[��������ӵ��FE��ű*��bD:��JwJQ���`֜y<K[����]�YT<`���lC�o�æC0�˫#c�P'�� �M�&���c��(L��,���)97��H�4�R��5��ҭ�*"�ln&[�����ޔ��mXRˇa3�z>z��ǋ�QW� ���U���k!2;S����ʫ�uq4I�8XKs�VBR��������NY����{´@�ڥ�$�6�Ⱌm���O�K�6���qa���KO�ԓ9��(���W�G�Ὰ��;z�tTuM�c�����U��{�y-���::�r9�V�T���DQ�rb����h�4r����俤�˜�1�-����(�J+<�����+j��kau�|�1���E� �|�l�݃8Bpi~����Fзh���f���NV�\�鳹`΋a�t��J�v�<t�jT;��b��*�>Ó��&�u8�0�����l�5��:�ZPR���;��g��PXĦ����4����8�͏`X�Sf_��� S3_�B2���"(X���U{÷��aso��WbC�|�|��rRL ��ψs�:Ja���eH��OS�׿��Sƞѱ�K�hd�&��yY��a��a��=^��(��t��	S�/�G��-b���>Ό~,v��P4�&���z\�^F��l���N�	����u[K�g<Kmt������]�[����` �ڒG���B'���c�@9�(����J�WCn>�]�6�&?C�U0�+�xL/����4TI�^����Ѽ��U�ʍ��M�.|ԗ��W�Z��#9G�#	Qt����0��v2�A�ϧP�k%�wE��*��cQ@��0��6?q"�����H��}H�8��E;�R}lq,=�5�~j���9_X�#5Lȋ�V�z�-�ba\z9vwu�(�	q�z��yu��1���9f%��v����1���K�JTM��%����TߟI�Ev�PwD���YMlWR�>�:���g�L��T�-4�ПP��c'b���͇�?]���_��ٍ�fIY�D�U��ە{��F�Q�)B�TvU�2H��r@>�h',@\>�0�ҏ�A���솧����Y�[�%h?3িR�F�	1�Ct��(�)����`VJ���l�oi�����٫Za�hW��|��y�0v��>(�mmƈ��tW�
�lw|�JV�E7�_���H��5�٤�:ܘd�Xc^�SX}�9��"��|��L�y:[�YeOq�)��w��$���ޖ*U~����|��O��2�y��J�In"
é�
T��Ź���)W��=��;��"�Cb� wo��ߞ�K>fO�Kb�I�+ʊ#bզ��1����F��!�L�'���^�?!2��e�Dm���;���A��ю@�(�n��ˠ&(��ket_�/H���h����@Uu����C�t!�5��6���Ɲ��Ii�u�D$"�����щ���={AiH��Ǎ�������:��
�9	��.*�i{L��F�;�t�rc�*еI��/��Mêl�
�z��)�ת���4i�~�����3$�O��#��afylZ��P����������Eq�,�m���k*��(�=qW#Z�F����
�aY�����zX5Ѿ�42aؒ�Iu��
Ξ�lġ@��u�qZ�Lќ���V����D�򊂷<�֔3��r��,Ĝ=�&홻�;?��V���f7NHP5��7�� �ex�lr���䆳��<IR�v���� g��b�$���$�ho�D�V2G=q}�
�T��BC4�ݒ�F�\��t%��O�߀�+a������gL|>
����eN�LX������&o �#�NC�ѧ�p=l��KIZ9�����~HN\*�qd��hB��=���ͷB�f��K�O�DϪb��e.�e0"�60�X��m�*��N_���cpE��Xql$��5���}�+O�f�[������3�S��1Ӳ�bB��ڪ���w|�dj����j`��3�:��s�4{%Xz�q?�/�ޤ��ct����P�
��᠊�]h�\Z6�����9Zg��Ԡ)����7�ΤA�_M� �juv�Jn�R��fZ�t��O^�������k`> ����q����k���VC�_|�5Q�3��£�Ә�/Ԃ���@��6�ߪ$�^��)19��ByG�t?x]�8Au���V�9���b}p6T�%=pf����P 6�n�u���8�-p���cV����x��X��P�{IYo#��6*�.��d�����G�v�B�(��@_���{��۝b�sʹ*��Ӿ�ſ�v�J�:��s�ޘ��K�= ����M/�wc�,.�a��am�`����d�em??-�J���Ԩ�%$X�f-�@�	��}�d?��@fS�w����F�v�`���^q��e��Q�j�a��b����ݭ+�J�%X������f0�|�6��>�Y�rc��~�9p|ͨ�k��H�5������]-�D��>�����4��t�h�RܖIǋ������y�@ҩP������[�@��"S��I�}3��4�����	q� xN|�䵩�އuX�N/����яja���>��0M.g�%c<0'�����Na�}�c�~��Մ�	��H�*e�+Y;���t���p�f�g����)��Kq"�Q�i���P�|��= ��-��2�mE���
:�_y��uF 	_vy�˨���%��:�_� 
o%�c׾W�Z�&���F�ч���0��pҍ���e���#Y��zܡhl���'e���*b<k��G޶!���G�-v k�Tŵ�]�YR�#c���i$ӊl�A���=�����x��E��҉�+�JI�Y�$��'C�� �[J3m����_����F������3��v�L3�7O�A�Cgm����JXZ�s �v��W@�\.�p�U����"w�}�DA��.���j�;/ �-U)��q%�E���*"���k��<S�����*���&��5M`ڇ�D��t=���-��6&ˠp�n�
Sڨ`L�MteM���]_B�Z�9_���?y�㣯zw>*g
�-��~�il&�U��G<���FL����X`�V��0�s&���Et��|J6%�STҠ_� �>��Sc��Wb~������h4�ZG�M�+%W�t�z�'�#F�z�3c�[�1�MH9����������߷:&�s�Z�+-�P���UcKx=4������hՅ�8|��P!u=x,J)����R�K�E�9
����#�
��p�PS��ҷۘkFd����2��˱3��L�1���|����թ���%Ác�m~�;�8�Z���H�_(9�<�p�*X8и��V�r�sǵ�=	��Z�H��5�F�_eD�v�ʑw����;4#��*�����7f�4�9e;L�VG�z��}ïwԊ-�^e�-���yTQv1f�-..+F����N�U�)��H�8O�NӪ�8�CP���K�Yvj�p���r�(�7:��~ɥB��o��2m�Ւ��_��zjG���%Y�?�I��w��<��DU��d��	8]�ٵ��X4~��컼|c��~'�U�z:s��]2����X�����������"ǈ�����w�=�
7 �cG{��5�[.F�g�&��/C��f0������E�V��&��f�s)Y��҂�$��(�_�i��^}�Mt�K�m�<=���)9ޮD(��3�����[��"5�����5����#c�pm�e8:��d'蓝�z>A�S���;����L083����j,���]�pn�us1(I�2�l� �
z5|Ǽ�6�WfV&(��m�h�!�d�̖��XZ�0ï��V�aJ�c�	 #
�;��{�y0 CPj��CH���\_����5�O����lScɗ��8Z��+��T�z��
�*����t�5���)��+��h�슝Ń(:=�v���.��U[��a��H��$�e|���/��zU��O���^`�9����s�PJ:佀,ACr|麕���7b�����Ӊ���}u�-��e%�֕%��Ioy��d#�qڐ�1��L(׊d��nrF�D9o �'GH����d.��ꘝǡ0�j��߾������4c1�, ����H��tѿ�S��ýf�"��M��ڍ�[���E�P��l��6�H��a��u��N޷ZN?"ƙ|=ʲ��}*�~.Z���jc�(R� aY�^�
`�(��U�<@tc��_�0�-��[8R*�����PW��X~�k���<!1㎵��i�leŴ�z�l��!ǗmKZ�!��)gJ�JJ2^��-/�{� �q`2W���K�5��w��cQ�Nr��=���j��=U�j��T0�����i|����w��D���m����狕 '��T����(��l(����4���1����y��\}7>!<��G����_��i֞�<X�o��aR�C
�.3��[Z8y�R\4���!s��r/bF�G2`Y�ԛ[%��8VpD|�	�V8��Ϸ�>���^�����[KpU�d��"���&8p�� ����!�|6$+���)0�)�^��c��YAZZm� �5h� ��ɖ�|���\?����������ZDRvA����^0���f�I��ph���0w�B�ҏ���������'��6�y��'����������l��{	�p���Ӱ�KN�||��Oz�Y�b�6 �@?�x�:�+������~?|���U��zk��ȻZ�����`oAH5��TE=
е�����P�'�£7lO�#��U��vb=ϐ, ⾾�g��2������"M�����1#��W �A�������"%f1 �@��(�{�{r�c]_�aݎb&���Fs��5'�u(;�)�ێ�Kg��e�)�:"beX���<(�� vfL,�i��H-9C�H�;�|�",�{��89�}zӎ��ҋ����e���c=3+��S";��
-�&�gn�-���*��"gS�J,�`��A�gD�i�c�5Q���C�	��L<K�@j�Q���SQLa���	���P�D����Dg���&�ª�jl�)���J��+2ܫ~�R����s��KS�! �$�@~C�Rf��:�;��Ev��S{��%�QA� yX9�t�U�;p��%&
�.�F(��>i��*���Ưd����L\9�}G���X�<3����S�����1���0�1��42S�9c��g��bmt��hBԮ��jS�o��%��[G����Z�tܲ�Br�/+E�=
Y/���0t=e1�:DfJd��/�Z��p*�4��˓2��޺��oʯ��-�E��
>�y!�$aiļ�A��m8/�U�+��_`*T�Xii���g����!�D=ɐ�&+����G�ж��9B�{�D��!�6��4��lQy��&���s���7	50s� `�p�h|�yع?�r9�i��RR��3�Y�5���pm���3���c��s��nM#0$����c���?V�=2vt�}޶��de��}�N��}J�� �F W��x�Y��\�Jh\�G9��\|W�=c:3�
���g������t�=��g�0���(E��}�x���p���U?4�dS��o�'j��h-]!���N �(/4��}:���`D�0� l�Y҅��ON���|jb��������i���� 0�X��뿬��%���e8��$�/C�tŒK��^PC����Ȱ��R�B%����L_���Qj_��4�V:
���;�Qiw�o8���X��\v��M0_=j������I�G5�z� аg����=�j���>)��ܥw�v-�Z�-[w�>��턻�}��.J������M6��o��u���[�\�ٓ���ɸ{}_Eb��uJSX~���| t�Ę��S@�����w�̉��Bw�z�Drt��M��/���p��5N��?	
byD��0\�e��- .!�2��TG���J�R@�{�l������j|�����9����_�mk;�\�p�:�b·q"1:�4�W�|�i��@tƊ��:O��l�h�%N����p��+;���1�E�?xeZ��aÀ��*m�,:��I�h�  J�c��HR7�} �p���
%�1�~FMŦ�P��C]k�@!bp�a�|Ig��EB#��k�㙙��2� 	C���T��s������(��r���n_�R@;F�*ws�2�PF�e�s�ʥ�����U/;���ұ�����2���UY��S7]m���E?[���R�I�>�_	��J�(ϡk/������	+��?u-}�<L��e7��sM����z�h�'�{�Xˤ@?����#���*�O�v���z#̆��ڝ����Qd(D�iq��
����?�3���.�2��L؆R�/[4�F��6�{����p6`� 8�s�q�y�{�66���O�ɦ.��Y6�P]�8,�Q�^��/Ŋڼ�W�'�ajQ�i����+� ���V���_wG���θEvnFqA�-�A�F}j_-۳F"�Y�FM�À.�Y��e��8t3�X8c��~��7#��j<o�!���<P��̱%�\���@�AC<ڷ�-�v��
)W3��ڰ�a��h9�����UT]��jpd2!�$�%��%q�;kz� �k�xEv���ƕC���q=� U��ىM%מ�'�=S�]�7�Cq�������� y$(UƧ���GZ0l�P�\1;�^�)2G7��wS�`��E�/�O��u�����zO��<:�z`0KȧTf�ۢ�ޙ��9�URgʊg,���ѣ:k����i�Њ�X<�W�T��lr�QaG\a �pسˇľ�R������c��(�[���C6�ҁ�Z�X��Z��+�@�84�%�pu�C�Q��r2�?#�h�����iHQU-E43:����<h%�)'��Dڄ�3�ʟ�2���EC��3C��d�T`v��R�V�P&�[�-3�L](�}:k<=��������A_�\�/.E��VZ1�Hc�D>�-�gHFv/�4����u�-8�n�ñ����'�k�� �	�������� 3e��)����| �'*{������sv�]_'�z��������]��*��#��i�0����o��L�:�B��m�&nC#�$��0��S�6�n�6n4�`�?]��p/�g��H��k4eo��cYք_*�� X�P��Z�W\�H������!�դO4�YZ �rϾQ����c�Q���P+���|B����\x�c�]�e8�R�A��}����2.�PP��<u�� ol��ߠS>�N~s6u�1�!s��9�[�n��ȭ�i���+���(�V��|%��1����zX�$R���kF� N�پ�����B	T~�� ��cB�
*�$֜�a�ZD������ۣ&K�."�������*��ѽ���a�1f��I�a�M�N	҃��C�5sq�y}h,�kG���I��h��!䶥�ʅ�J�f�#_Ŀ~g�WBd���E�b�2S��vJbY�rޥ�[�H(����
��&�7��1�>���6n�ޜ��pe�/�/�@�@"����a�ߵ��d�;(����e�bA��9d�7(��Y���2��JƛvT��5��n��At�zZ�R��)k�@֗���c{�A`��i�d6���k3�%���Ƙ�>�^I�8nL���O���N�R: ����6\F�W�N����U?�I ��k
����9�%���rư�<I�@�r����V]�G���{5*�p���M�}��(��s�6�j�:*he	�SibǺn����*&�>�܎[!qcLpL�Đi
�Br���s� ,�P�F{�S>�T��=54�A��<���@��U�'��dJ�ѱ�k�D1x�T�<���'o���ё[�v�!� Oh�9S"�S�GW2EG�|���&b ��3��}o�u���x7��TR�a"oWv�_	���{�|�����8���������x���E��0F��(sA�� �#�R�Ȋ�����t���7�T�v��zg#�����'�����q�[�9)�܅nn�JXSV���`��i�B6�r Rv}�pw�=n�?*�܇66��w�(~26Hy�v�e��6k�X�|U,ʹpN;�95�		�D#?MĊ�E�=PZ)b΋ec��NiDx �i���Wpok�7_k���k�{��ș8&@���C_����
q��f�!'�.-�Ǫ+�L򥴒L��݁��r켧`�#8�C�>&�V�[%T�G��ԩ���9&�D�A*���њ�\$z�#���X�\8�ɐu{�'^)k���8��J���>��y�;6Ӱ�fmo��Mp�� �e�PV����� ge@�K��ɲ)"@ l��b��ݬ�2�hi�8"���R���-p�
Z

�ג�
����#�u���`�,�$�[��K��ǅ�8�ݯ�럕�l���i�|{,c�
�V���i� �i��=Sț�x�4��ú���:�����xqÆl����@ou��8���KzEu*Te��(T�I6��I(�f���2��WB��c�m�Ė�mĪ`X@T$�W`:���������w>b95@���a�h~h|pz�ۆ�	���'2�1�F��~)�r��+I>#�Ny�� ��Pu�|�<��vŕ�0js��0���_ހO�,@ߠ�Wm�X�GRB5J�X%eIUxM<D��b7���B�%�.]5�Z&��=~F����$ Ű�jz�:������D`*&���������p�Re�ݫ�tm�M��;p(��i������6�n@LYC�@дd�Y�W����7�I������~5_������-C^%�9����3��N��X%���(]zӅ�����a��*�qj�ƅ��+yT��w�/g�q7 ๳�~d�".lmA&��h ^k*pI�1�چE7s���P4ǖGGg��������e��r}�2�.�灗�2\�<�SH���wK�W�W�r��)Dg��XI�*u���P/�`؄]���u���ۖ'6oJ��t�iu���V�R���!_N������fPSz�5���Z��3c���X+'3I�ת�B�G��p2�=�Z��ZT�>��а�����nQY�|���� �{5Y��gWq�s�G@���t��i!K��V�.�� �g���K�>���X�R�f�H���&��/�����87�'�p��V,�q�frJ��td�����+S����0�1�Y[3�KLQ��ȀV��ZI�5�-:��/���~��4�>y�I�\�ilQW+������d��2�խ}�03�IMf_	Q�;��*ם!.��k&P\�\�.m�h��i����աV �0�%)��YǄ��t�$�ۼ��	d� ����^��� M�55�3`�8� �DZ�p��{���Tϯu��PrU�}fx6r�qrr�pf���Y:��9�Wd=��*�77�=�k�J�nj: ��Ƅ6�/�@���ݒ��Tñ��%�k�U�b���q׾��(�����0��j������{.Fֿ�E1&����O���Ƀb�t>�0s����#�#��?�C[��Fs6t{��7�f�7:\W��{c3R=�rs��B;>���-Kd�ً�Ӓz�+�DD@��OC��0H�����~�C������,zw��%�90EdZ@\I��B����;
6�Jۓx���<�7����>l��MG���I���W�0�M�مk�����}�*�ތ�S:���ɺ�1V���Y�C)q9�nɘ$We�4�d�X>4��M!6����zo��՟�B<\�k	WgN��P�7�!"�7_���W�7䥁����+�
"���u����E�[Đ�p,m�=-�K���㲫�Ø����u�̤y&TL4p`�a��A̨����z���C��?ъe���ח8�u�]�m%�O���`��љ�{�t.~�W{ y8��!K�C��1��݃O��Ș�Ы8�)޻���M��%��lHn��m�ʥ��孿���䲪��5�9��sv�)ۺ�[�����;7�]��룍l¶���3���ֹg7��?3�֏��CD�<��~�Ӏ�o�@y��\���ʖ�!��!��*��X!�=��{R*d&D�҆iK8$O~��-tR�9�i��>�z�3d�:]H)�~{�F���K��T�οD�5zle�ݸL����*�(�@l�٪5!W��YUř�Q�|?G����Gѻ�a=�қ�Qde<�&��k��P�L<3�g�(Y���2��M��7�W�����b�sg�G�g ��P1u�7��8�p�%һ����;�0���R��tyX1���;$���B���!��z���<�	9��"��AR�S-5m|1���W ܽ�M
�adP������\�ޑv۴�1���Aӿ߷���Y���Vcf�oq�#��x�V:��3�����w��Ե�H�f�$_����KA�M%��g��ZkUDdP����U�>=�\%������\���9�͏�x���϶ߨ�I�L6�K�"�ngf>��Kޚ�����Z8�SQ����_C+A@m%��-&h����]���F�ysB7y��(��^J1]o�v���H�D׃�d������ S2��RvHn/^U
��@Q���faKZ6R�O)[�mh*��UJY�D�|�,/]�a^������2X%�QM��������=3Ĉ�VR�=	{�}���oI�]�Z,η����RI+��3|q��0�Ff��T��ꩈ�O��)&��#a��4�S�U�v�Ǡ�~��� �3;W��0��S.D㠜>��ആ �E/�����λ]U�G��k���x�ݝ�i3L���=�����B?JIEE�p�"<9��HP�h��������,�0*�ߴ�D��%��� � [�<�o��k1�К�V���{��/@�x�hN�?��r3ב�.d�[�����F�jtPq@�� ��뱅��u�;R%��������i��u�Ŕt+�]���%���P��'i4�W�j�uD�@������`�������D��n֣t���a�"5Z�i���L�oT/��\KI��NßHa?�Z�y8ej�r����u����!֌)�q_��W]��}�h-k���P��a3a�S<�.�:8Ҡ��% ]ta:#c^�v�Xp�j��p���j����E�X���=lq�g]�=+M���f�ۈ愌zwf��1�#X>s���p��Q.p�`4�����a�(��>��F#�3� ��T5v
�V���/���)�ܵ�V^����Ӛz�*��r�+#�PYJ�G�-0Yzy�Є>�%��;=#5�ϗZ�n�~�N��+	r�4y�v+Z��ΥKW��Tm���a$� 6�k��k�f�V:5�3��'~	d��dA�( �˂ߵ�1'k ���x\�S�崆�e�����8W�����zp���}|V�L��b,����� n��(	A��i��b�̜"��_pД� ��/�l�K�0����$Q�:��+!��
���7*V��k��1�vC�u�L��<9�qa�j�5�O���D�N���Tik��~�WA\�0�}�\k�pQm�-�Fuq��kB�͏#s��V���bF{�����26�20y$01x��q�7�ILL���I��[��mB*Vϸq0;�0�E�q�E�"��@/
����XC��L��=;EJ�j�V��p�2r2� �@� ˩����O/���s(>
�.�:�4����-gCP��kN�����=���g�ʯ��6Z��n�����9_>��ᨠ�?&��K2}��ܩ��<nŇ�ԓR��x�H|!��W� �̅��y�p����<c5�s��^��[��wAx*��Ī��,��T���f�X[j�2|�V"$�9���E���������)i��*������`���6렌`��s������7^v�:i�e��!�(�/Cx�o�`h��b�5����?X�{�_3�6����^���hкb�x��+���z$$����K�4��5�h��0	6�9�R.{�F.���'�<�'�iT��c,�*�/|C��h;lE�Mm|�}APD��6�ϑ�V.G"���Om2=J�K8��������>g8����Lx--Ӥ�1�;p�{e����js�J���L�-�R�rH�8���v����-�J��;0��/�h�S�&r	8bC�l�Ǎm2��vaI���mM�V��e�Z�b\�.Ș�g6�����I�Z�AO���oT�Uk0(���US�� =��33�ǒQ��S߼rxe�*x�~PQj��&��E�T<�
")G�¸w�2��x���+���t��ԥ��p*�C����8�3��&*w$�"�VŒ�w|Ԓ���b>'�_�C�� Ma��w�tP�L` j����&�5"��V�}cEN¨3��70�� ��q��X���$|��c� $��܆$.�(Zr$P.���>��Bn�N�/��7䠚��T�E!m�A��k[ƺa;�%�g�K�4����| )�%�����B�����~�f9�-gG�bbK�Ut�����Q�Rn�F���G��t�6K3��[��z���}��f:�G��0�}
o�0���`�Z�C�%a�R�E��ڧ�pP�$�'^
���<�?fR��ؖ�6��C����X�
H'��޼�rS_������9B_�a�J��(&�Su�y$$7灤��'�5��w�(��sVxhb��roB�bw�Ps��ؽ	?.���pZ�=e6���8果�Bއ8�����w
F�6��?],��8,��S�B�a"n�7n�?��ݲ�PR�g.TS!-A(wj�� D��i�-8���IG�؁fg}������C�����ґ�ߵcxi�.��mE�	�c�p�q�Rf�ְ����&Ujv�]�����������6�I �ez��x=�/�8�!1ݒwm�93�u-�,Y��ƹ�dfK T����*��՘-�CI���0��>��JѾ3S��
�^+��ris	��Yj;�Հ��Z���{3ط�ȑ�����6Q`�<?�Q�C]��cKS�k�0�i�L6���zM,���؛?#�2����8<�]���v�|&��D=i��&p�J?|����o0M7ʏ�#��KKv���W�T�WB��Ox-}]
wҏ>�t.��n-���>4�����/�_�^�ׂ~����=@ �0��v R�U'FD���|s�J'/�mw+�W���g�PO)2.�N���h�'q��{��S�k�Ҍv;�O��wx?�����SLfX\�EϹE��Y��<3�e���N�g���f��90k*�}:X+xŊ{��ǰ���P�GG�����%[YB�O�ps'xo^A���O�qg�6�������+��T@AןU����l�:�cP��cY�=֯G�e����?�`=8�Y�s?m	�t��UR��ˌ��OC8NȔ>�t�r�K��i��%��4�
��e����(�"YX����ۋ&y�4L_o�����6j������DN��]���	���~R@��J��g~�V�1�����+��9쁋�?ڗ�����.,�!�*��S�rO��7�� Ѽ�9�Y��B�Zʇ�6tL02=s�Ma�M�RG��i��DO	�P���5��~��O�q��ڃ��@��
s���ތ<��h3��� ��v��0�Ë���s%�ӳ�ę+[+�n�!T�sW�S?�x��<F��̗�<x�Q�074����D���������L)�?ko~*1=�&{4E䢱4���9��ɍ�8 ^�#�U`ï뒏~�󚣺,zZ��,�����\GU)�,�ll[Y0��p<�j��2̱HᗓH߮�hM����N4����v�&k�_��t�]_/��C]N!��Q��o����$`"@&�ٕ��G��K@�ѐ�rR��~fP}��ᮯ��G��J�!3$+���ַ��{4���11Z2���n�O�yj@�!��Ckc5w۽���;0��2M~Ғ�aR�,9"�	��^���A!%�8����F6�*���ޙh��R��w�M�R�5V�K$�l�V� ��U�`�D��yP3�6�r�x�Q��"�̞�#�{��ok�߄�Ʀ��/�h�YY�Sψ��A�	T�`#"�S�Vj��@:xi��\s1�~�ʍS�e�}%%}�Q����^�>�$����$.���q���4��ǂ�S�ϋ&��wAlRr����=�֏���؊�o�����¹���G���R��8Yҝ,+��A�q��_�`���4���+��'��QC^g�K�gn���P��K����Ӝ��_ZFg'��m�`f�]+��~_���pζa�ӫ������Q�U���Lإ�6��'7���sg���|�!ȃ�+A��\9}�:6����>ڴ�[W�>�+��)��J}DZ�w�⤞Qs�8��:7݂g���?{�Y��e]�����ם�������r��(q���~�a��v)�IR�QP�q���QAU�C�2�i�)���u��x�##�����;������	�J)��*'3� ���3q��
�@bD@�lw���=���O���)�&����}�]^�n�Hm��w����Dg�7���U����z�@��	�r�%Ny2G�'�,�s��G�k��SCi��iF��Z'9[��Hks�A ��ĺ��U'���ճ c�ѭ0�$:y�:Ћ�'�/�q!����k�W�eWnT�{���U��A��A�39W��>}uI���L�5R��&�-Ea��ƕ4\���v.�>ڴ��+�p00*4�<�.�ݢ��@ʵ�����Y'�TD�5�l�FᘢY3Y���.[z���^��\�`R�RZV�]ҏS�7==3���Y�]�y����w0�&�<��]m��'���B5�G��6��*��ЇV�I�7�{NN,���\52�X��ED�<�*f��I'F	"��vFKF��"����ej�����d���s���U�>���L�; 2W��"w"���e+�B��wNP��%]ע,�l�b�N�%V�#K�Gr���@�!����U����זu���(��"6��(q�A�=�o�6������N�E/��^��q�m��\�a��`�U���#Z�ou��1Y����';0�t�C�ɱJ�G����G�4��� ��2���*1�ӭɢ�x#�>.ɻ5��um"a�O��� _>&����>�	g�I���B�'�;���v�6��.����W}����q`�y1	�*'�E�E���&�oϢ{��u����4O�DV�Р�E�ڿ{W$�>�F�ܹ7n-�������8
+n�c�2�Cu��Y8�9���|�2J��_]�fM`' M�{*����-�{�t�h2�o�h�n�d1"ol(��#�+�;V��F~V]rPO�ߗdnjg�
%yxޥV}�r_�a��:�p��a�(�Q�0K��:OC�kU"�,�YU�&-TD	��a��qH�d}�,�ea��,wH��C��s^�e�?E�[��0ǀL��VZ���y%����z�e:�����$�Ń�m��������W�H�����\")8}�A �ժ@ß/�u�>!�Ȧ�BwVk�����YL�.��p�v�6�g۱g���"vC�'P:8�z}�e�|����h~����}�O�!�PeC��wЃ��f5�8�XS���G<L���8�����^f����/!�6�m�6<�S�H$����om�"���#�o����{�x,ۍb�0 t��p��
|8�tGk��o
�oĲ��
�{��
�F�f��[Y�Z�Z����|��0V@#�y`�@����ĵ��󟒜��c׵���ş��}���2��&�]6oo�[B����1�?��.=L;�8u�Fo���8�� ��oL�*;̒n�V�-�o6󚺑�������dfXX�(B��P�+�R�C���D��O���!ј|J*#OV�f1'pA��7���W9� bg�8��-�z�IJ�IX���j���ݖD�<�<�Лַ�ɩ6`{>f,��f�� F$[�p��Dn�XY��2ًTh��؉�=�^d�&�6~�B����xW�7Jb��L�!i1ʯ��&���뀨S_({F��ZlL�����.@�=
Z��'�[���>�]2�0�+����M~l�f�;�V�e:])����b�ަ��t��MK�ӽS�*qbŀ�\l������k��P��5Q�|s��O)�l��wb��$�a�j47�	��(ړ/o��,K%�!B�:�F5L�݁�F��� $�ϚI7<�_6�q�ԍ���\5������³vF�˪�
��Y��%aeX6Շ	�O��.C/��gR��U ��U,'�͠/Fc@���`dE�.���O#����Ain����ĥG��V�x�pÞ��6k�L��(��sJ�����}�H81]&hYSط�яR�����'��.��X�-vd��ԲVc�-�j�C�۞�9�DY�쫐�'I��>�c�A��{���F���p�"�d���7���ee>v���Y�'��$q��n7����B��r�I�ԍ焉?��=�5Ai~Н�e�H	48���O����$�R᧸)�q=zd8Uv��*�d�'�4D'��
��`VN���_ը�,,A.�"#Q���x&�&;%�������4'U����I�yL�)��k�������U����y�T�^�W�e� �P_�{gD�Ovs�����t�X�9C���rrs` N��� ���������<9�@Z��k~�╻:�"�u�}?T��t/��V�-�����S�i�j��7WL_�2��k2�Dփ7	l�q�L� �=�͗eFЈ�_��j�n�Z��,�#� ϱ�-l�A��*J��{�<���~�����'�d���
y~���c6���g�
T����5(�<�\�A�#��﷢���(O�@܁�S��7`N(u8��e���?�C��r\Q�(W�ٶ/�&���H�����#˷.\0�o*��<ۄ~L�
���k �vw��K�t�?�l�vk��
���y�<-����w����#�crq��z�:���^X�(�Ǹ�c�\w�����3��_\�D7�b�K��4-�v~�����_I_/{H�U\G��A�<*� �^f[�)3h؆ u����C!���g`'2GP����4�=�C0� ����{г/�/�����ӣG��nY*�ˀY
ȁ�6%���`G�KRe�a�G�kd=� �2��9��r�}�[�O�0�����N3n �J3�f�<�<:@/���7;!���]��p�yCF�V-n3�����{����"��@LCg-��[�9�@�p⩹En@3+'��Nc�33��t{�A9�f�`��$f���b��8 ���f���E̴V4>I�����.�����C� ����A��ε�XHs�zC���ԁJ~��<�Y�1�Dz�lOK�\*��tA#���5"Q����lTdqR�����L�/�j7��7��y�訲y�ؽ�%�Q��Rq➂u��Y��  <K�E\�vX�āK���f革��t>Az�?�j:�Y��9�N�¯U�m���"��oU~n���ZR+ĵ t#P|	�:hxэ����f�*�z"�w�`+5;<S��d�6�����)���F�6�^�A�Qo�y���㏗�mj����;�@\_�䵟���&y�Nk&��^>ψ�ȕ�k���a��:�T��l&��@R�ۺ��7�<U)��m*�L>����,��lnz5��\HN����HIT��"/����h��ٷ������A�Ȼ�a~V��9����:Ɔ��whN���t�C:w4\�A�����RM�]�������X�� �*�ݓlV)I<��m ����C/�i�A��J`�2yS��gP"��$�X��z���BʭSkZ��<��V��VZ�@�9�rC>7FсZ�j5��&D��Ӏ-�l�t\ʃߜ����F��d��/"]���<	��IxL���1	@�<���	p�,���$Vֈ@��	��O��1qN�<���F�5pWDt
���f�F����ey6��K��E���[o��@v��%�kҪ?L4�N�;s�#3IZ1Z!=\���,ІuN(��W�/��$��]�~�eڠ$�:�=@sup9^%����!ْt-o����j�f�E	.��J(� �?����ݲ�,�Z�b�b�n�M%I��斡P�0�Z���(~q�Ul�{�n��q�7[�a��2�6?�%	�(">�����ј\x:��3Wdd1ˡ�<Ԧy\�7�3n�	��Y�<�{K@�(��iI��-و=����{� $�Xl*t�폿B����.'�S%��5������xi��m	$�@�nko!mC2�.���p幆RIǛG��3�=q����f�(���"(���!m\Kd2}YK�S�J������U������7��\/R�c�icx�	�9��SƳ��+�!(�%���^���Dl=����?���H��up���%i���+��& u4��,�	�h�/i�.�o�qɫ�C�H�\�֬��u7�"A��!��j�"k�G�Z#m�Ns�d�M��X�5����qag^��ǤI��d�>K�Eߔ�d�Xuh�	�,�%�ėS%b���L�TIXe���Xd�o�\LP@
a���!��:�'�ǅ��稪�?��0�}Q7�u�V�m'�x�r�V����e��&�_~�K?��P��� -�6c���!��C����l�$*<�]�c�C��Foؼf�aņβņ��"Y/ ��Bs�`cYc�(�2��:���������8�̀�X��A^Iч�L��w۬i��Z�����Z��"Q_c��h��[�k�߅:�K0 ��(�W{���f�|������;�w.�����Z$�\d�OJ4�o�A�l�p��>'v c8��e>����(g�B���ˌ���3���\��`L��� @BY:�ّňpP�=�z$��Zٻ������J|�����:Z� Y� �8��gJ3`}Q���겝Aid�X��e�=�v�e�Ы�� �qR䊲\x��a�y��a��qWt�O���&�W����'��	�:�s��jɥ�`����'�v���i��oF�q$,��4�M��͟�	���7����e� ���EF��zQd8쯈�o��Iʫ9c�D4�r;ƢY�a�s+d����UC���9fwN;�hCƺ��S"�4[s(
�-�+w���F=ojqzȮ�Zk[�����Nn۟ab��e
��S�b�:����r���2���֠�}m��~oo�>c6���0z21�p�Z��Ψo��Jz;6����-2�����$b��WHe+ɧ����{>n�N�O����j�n,�F��p�� l����b��-]���?��Lg�v͂�W�m5��G,�uks&���ː#G�J�]���.nռ狶��*?y�\�x'�P<ƙ� �JNSl&bs��CBeIj)���I�����9b%���3�`ґ�qX�=�-{ q�'�BN�@������[�=�ֱ�X�#���'B�������p.?�>��~�ΩCg/�w��[�y��:A�0�HR�ɰ�a:n)��:=�Tv~��`��\i�K�alz�S��S�Ly}��)�0��I�q��xSeQ?1Sу�9b��߮p�}�.�b�	��Sˌ�7r�qw�	�e��Y�V>�5��<x��D {���$�卒Bi+����el��!Cy(#�p�vFn�M�.�$�r\�^��"�%826� �|�C�Z{��z�@{5�C�E���Л��*<�p��4�W���5��~�l[&D!c�Һ̭}~1�O�Q.3���0�g���+pi�+	rK�-"�ckky"��)�Ak@���N��DsN�4j�ജ����F�u���� ꌬ��q����3�������v5�$��ZemݙR��T���U��{�Szh����ӿi/|tc�܅d�ga�L���^s�4���z���zp�Y������{��
�YO��I�Ee넔%�_m��M�d�";		'��Nv�;��#�lC�׳(�M�<�� j䟮��"���C�oB�w#&�e]���0���Th�i+�V�S���F��[X��eS��6�%(?��s�۔4n�=����G2��6����
�3�9ay)���:4h�:;�z��������r�[��X����{�HMZ���b�[��Pf��.O�5K	�0��;�M-�ִ�\K��l����O�eo��3�s�<�KG��H���+8w��~��͵n�Mt�G4�p�r�N�������pn�w0�T(N��n!;Dc4ysR!w����l w�F�>\^&�5w(M�rp�͌dF?$���YsU�7F�r&��g�L=�d�-S���Ʋd���F��A�[҇��GK��OU�4�H���l5(f4��9��{٘��'%�� ��%���%T!B�*����� �DmPF��jq�k��J3��Y1zԣo���u2�8'�m:`5��zZ%�ɛ�:����-S44tD3�~���_@�(��_ÃhnJ�^����x�>��^��zD5�1X�z\�-�3-�B�uW��k/d�aCX������m�ss���<��-����z���D�C_UL�JK+A�{ۑ�8N-���͓�b(")ѿg~��X
}䩳�S"\�`�Y�Cm�8y^�)+
� ���Z�V!�i�%s�\sg�e�9���a��z���e"�^מ09FO$�x���̭��s�]�,1�Bu�n�Ʃ���t[�T�/oS�c^��� ����)��P����7�j�"h���u�$.\�^��@XB��������	�/�ڋ(�iT�����1CT]?�h]�<9�����皉sHJ�W��(���z��쫪ڻtU�8J:�Jq�W�<���f���] O�l���uc>��)�B����8�O+L��d�S:ޮ���T�'�pB�Pm =��ޮ��-#�I���ᘋ�^�@N8-h�à�~�/��uJ��!�blŐ�п([É�A8nwEI�^z�H&�t�`pX�X���}�G�����t�+Q����Ɍ���%��`���Qn���j�����ħU��|�xƮ������}v��f�k�1A�~�C�LXK0�� �f!����L��%�A��S��U�sJNĜ���F�[Wl�JfT8�G�!͢()�#��+]�����{��e(Gl,��l��V�^�	Ou�z�� haz�W���&l'Υc���G���2�!�
�9���6N����:������ p�dPJ��l�ں4,����ֈK��ml�eHk����Þ�����"�K�U��t���חJW�1��$���,�VK$@L_�ӝE�^���qwT*Щ�|ieN9��=�S�8"�m��ScP'_I�jT*	�)$�S��#���D��}јhcX~��o��5�����]���H���#b�*��{�ÖϤb�u��?'	�A�pWbl�G�Q��o��;҅"�X�J:cFjO%�|2���dQty�h�7w߱ry](Tj~˱|�Um��z̀��U?��� �y����w��6���%s�g\{���o���R�,��pE=҄^.���_��l�
�eV>�K�)&�y�3�_�*��?KQ�D���l�꿼?�d4z�o77�>�o*�ӆ��y��)e�{<�H�\l�U�/r�������_3y=��d�Bp����A3E�2��9]�ө� ��pHW,�g�e�{BE�&|D��*nQ������D:BlB5�B��f��GF�;?NA���^@^ �4-Om
�O?���m�*���+X�-�φ��/�Y��q����s��I �B��-,�K�P����F��58��6N�5w7�U��YZ�2R� ��,�&&!�MC�1~�+��E�AT%W0�����`����Ҡf����๖ܣ=r7�X9��6�{�L�4���,�撂��\�zt��	�x���ֶ�֣j!:�S����0+J�Չz�j���!�Tо�ø�K�f[�8٭�O��"դ�U*�m�D@?��G�_0�>InZv���iS����p*tI���Imv���Ԓ��ҩ&-�M�e��FȜ�3|�TunO��q�sc�H��ٔ����Y���X��!���C��2��\=�f�P^@��-�02�,t%�Xg�T(�2�NuZ��V{=��8 `<G�b��t�OkY���i3�%���W�Yi�� �W�3��}]ݺ�F�~U�lIF�qea΃8�V�����z_-�Ua���J��$^|�a�/����4�*�]4&��^s�� pm��̓~�E�Y�шK�,h����4��*���4�8�'�'��@�1��卟bkk��(x�����b1�u�O�62�A�Fq�)�<��P4�2�����K�VQż�
����d�U�d�5��;�O�L�H#Z�#6^
5��_���10���w��#��S&���G���.w"-�L����Jw�{LL���a�#��H��?㋶Y*`F� X�.=�u�+�G�(��N��l���Nuԧ�kV\�Q�z����H�3����9��~��YΖGt.uH�L��Rɴ7�
�)� �Ѭ��3����A���T�io��Uj�lF�Hs�nf�A/��U�*�k����7��6M�W�7��g4����Q`/�#nD�hm��i|-��\�:/���>r$YGР)�;�`0b��w��m
�I+M�Y	�}9e u��s�r|{�?�p�2��0x�'�nF��q���Q���wJ]Ƌ�k�+����,;�	�(Nѩ�{L֜�0B>q^AcZ�#����R�j�`���a�O2�⥑a����ʍ��C����:����� �rזu�
���le�AH{�un^EU2c��^ob�\���)]K��;q�w�������ΟmĶ)�9&PP����}�ׄ�e(��Ƭ����j훈�\�n;������M,�{2V�-�� �n5 89n��/c�x7N�:R३u�T���`��0w����Њd�|	�ۋ5���G�i����7I�d8\��?&�q�
����ɪ��0�UJS�ԫ�Û�sU����[��&�l y��I�q��{B��@ᨮ�ݠ�QFN���K|�1
��Э}��J��t�:5�lp�&N�"ñ�3R �߃����@U1(_�!U�.�$�Փڸ$�҃���!�ة�JM5���؏�����G+B��D1,>ͩ�\��ޑK�����I9���t�~�X�v�')8�R 9Lj��&{�XpbN� ѵ� �5�S�"�r����M<$36��0a����ȓ��vcz=��Y�QA�N6q7>�B�a���Xӵpm��x���*��$}�h�]�RB��������\��|�|�{�r����<�2}�':]ka7�ex��KD�4�*T�'TeU.�+�k�<'uT��C�حǾ��(e�L�M�������6�G��P��*P"[F9_(b� f��3��)���#��,�h20/��Z(t(�-�Q,|���7��������g,w�����g3�T�W$(�!��p	��O�pR�cR�@�8Y@�.'���|�_Yr��ێ -biF_�[@� ����ff�c��و�H�Z�\%o��)��{b�ɉ��c�`,�����:�@[`�܀��ٹU�]��ٲ�D���N��	�՟�Y��� ���`gL8(��+�P�7����/���j=+�R�V��ܵ�M�s�r�k��0�*Xpلi����(!���z���5#��u��?�ī��R��d�����A1�*~&����v�i�~M�����	`X�O� �d-bi�<�)�n���]LO�f5��Y��D�2�O�*�zm��<�{���� �mYH^��'Ƀy���QC����M�^�{�n�v+����{*|���a�٥�[��� �1hf�q�>�o�͍{����l��rD��̴J���f?�L��9��p&q ,��CI�����h�,d�Ʌ�XB8�9z�cNZX��S,tF��t^��>4�nQ���d�l�E���1�n��;��Lj���O|��	w�S!#�V}��"�*০���P+������H#��+�ڼg-��2��
�#����⹀�q�^�|��'��ܤ
ͥ�����ܝV�7Lf^tEvp���Q<��ܞ	͍[xP�"���Z��WI;�d��ު�����.�4��Jj�GF�ag�Q6�TН7�7��&s�Q�B=�#Nb�yg�`��� [��
�h�p��;(�dGVtׄ��Z�x�$X;���`�wJ��i1,\��t�p���w8�6^�@?�[4zn�����8��XQ$��x�̝-`�*�s)p7�E��2��.Mv�rE�q��$O>1��>���
�p&�ʦ�p�{+6)�	9O^-A4�O1t,�":���`a�8�,F{o\�xŜa9#}R��G��]�ϕ�G���ѹK�K*��Stf��1���Cɦ�#�'�WV����#�R�c��C2vӎ��,!��7�
S<���Uao��*V��ԫ�
���0�*��m�zS�J�z~��g��R�g�퀉	�-���n�P+_nE`5�=��r`a���5�ֹ���?U�����S��pJ'�n�gJt\Z{,E�d���P�K���ʂjy̸��j�P1�!�%&�?5�-�'o~Q��1�o9h����AKUj�R��7�޽��K�P�)�В �o�,L��G��{~���g����a������k��0_Ӿ����,:$��XW(3�8�N9-��RT	坻�]���"�������D��qf�u��&�&��{��$�jƓOa��rխ� �R�Wq���h1O�F�4��S�I��aH�9��	�ð���I�Q��a��op������b#�w�:ﳀ��O>:���s��B/��W<98	�
n���Z�������n6�,��x�%�UمtPO'�HZ,�.�̊,�FAwР��N�~6��l�~F����I�����eLa2G����8�M'��=�V�,x"8F����J��t3��Z�7��hB���s|�0E���I��l�j\���TR�F��2\���zz$���R��jj�<���i�c�}�{��[c9�i��j��'i�ݶ�S�C�~4��4�����P���(_|�������/����`%���K^�����3�d/#\�s�
3��ʦyyhr3x�}1�����Ks����eATY5�>���g(�V.]�֓'�/3<[aɏ�
Lp�{�S���Bd�	M��k���j����4�UKQ3�㧓�U`��$�9w�ҍ(8?G�cOg�u�5˲�G�"Wߘ?�td�X�W7Okw�c�8O*�8��a�;;0J��$�1��f{��Y��z��f5٦�d�m��T�{�DZId������F��폥U�w�2����'�<�'��E˝���K��&#"IqǼ�a���}w$Ȕ�7 E�;I��t`V�_���1ɜ��@�'���TE_T� ��ͧ1+�Ѫ��0�mO6��+�=�P�E�c��4��@4��Wp3ܧޕeт����@zfFC�����;��ѽ��[o�q�����b���Ҿ��Si�Q��F�l4�r�����Z�%%����/u���-�n^�/�p���^X�e�T^�aa׌k�@�[����6�b�9��L���D塭�(c�K�|ȣ|����a��rI�}�|� z&r�|��S�r�� ޗZ��%�٥o�-�~���S��srѱ�������71C{��̋�z�cr8��[��@&&��DZPI ?\��^�<#�=�}%eKg�q��{�ZrĬ{���b��H��5���xR����7��B6�z,��?<P�F�^B�1��r��a두��u|�j��Bcy�Дɢ�=���������,p~�Z�����ޏ�a���Â�L��O�I���d�{��͗$ K0�O�9�D�� :Jہ�'g�Bp�.�!K�syzi��tuy���H��/ɔ}��B`w���B��'5�G�Nܰ3@���EL-?JA ��k徼��_ퟁ2ڠ�з"�r����Y��6��'a@s��ٲQ:b����(n�(�a��x���[�@�!�����S�h�<��Z�.Y3wV�)S�s��vW��^�S�B�OlςX���M��T�u���B1��a0�!O5���'���f���yy-��0+�x�𫘆��o��q�.8��:;��y6�!%��1�П�i?�9;T����$R���(�
}ar~f�!q��8��f��Q�=�?t��\�а�#�K5uq�u��1�hˣa��6��#�e0Ep���G���c�tR#Đm�'Fp{�ZsV&��t���* ��1[P!U�cnv�u�o]���
'��e>�e2�<W�|����"������u4Tp�B{��P��.�s�`�S'l��҈X���/_/�hYKWVJ��p.q��G� �,Qt�I7��Gmm�����I0���ҽ_U�V�RdIS7����+f����?t��Z�M�^�p��z�����m����ɦ�b�:���+�τ��;�a�>���E֕���f���� ���@{%_�WY&y�{ˋ��&Ef�`�LIנ`>\�#��}r����Om��~}�d'��sMz������PW�����LS��ގBb*��?�7cbi܁tk���j��nb��È,.�!O�0����HH��؝�o�Cc�3x�/�,F��d�iOE���ۙ^w�Ql�Rbؾ���S�=O���Ǫ�c(�PW��9�.4�k ��\+��x�gj'�X��I�\n2^�����$O*���3��2��4���GIR]9�G����.�A�aՌ��#��=�Q��K�rX�2��E����};�|��Zo��2�g�D>�1�c�m���Uq$1�kפ�cē����q: Յ�]hf�O��A��g�\+������5�vĻ�"@|���7;�ڃcm�\ ����Q@C�2�����spD�g�Kec}:�Y����"T��r�8m��&��X��x9�E�/�_#���H�d��*�f.�0E=6���!6a��ZPWhc�@8֦Upr8
�9�R=�v���h([ñ��3<k���["ghV����FK�� Oc���b���v��w��vO��J������ �L�M�@q0>�W��'����6�WE"%�[f��#{����	���G��ə䞶</�PeE�+������yED��-�z��H� �p�$����\��7R��b��2�X��0LH��vkW�/��f	$f�H��n��Z!oo�w��d(؆��3��t3T���/��V��:�ڄި�~M���?�y]��fdc2P;�T�/�G�A"5�65�1����OA!���th�:F�v�K+�k��|��iշp�tNo8��ű���L�������ۋ_��� ��M�n�U`������~U��N�&�y��)K|h��gI�C�� �/o'�e��'C8���>@�o���
S���@F���,uŘi`K�p�!��0�`��ŉJ��A����H�V�R`�m!{il��'�)rl��:�
F�RN<s��.���������>��F�0��3�U�����$����Y�Y���*��b\;*�~�#Y%��['�H�X(6>�&��d�{�Z�|;�a�o�L����O2N�pobK�4�ي_�#Օ���2q�ƴ'#��+W�׼X��J2�(���n�bQ:��h�������Ы��'�4��9�S�M�"9���zҊVA���o�G#)�d�⏾$"�=p@��ri1P#V�~�m�4�_�XB.�ܤ���d�̼"�M?5�P}r_kf���e�x���K��Q�x��o<|���ʭ�N�V���m�{�z%�u���*#������\��yb<�5U�R���j���BdT�V�J�.}�����yf"��ԔTRq�}������WSn����t3��&:�����E�Hp~�XM95�z�հ��+P��������G?q@V��L��Zn��	"Mz�zQ��΃|��M�j�E$y�;x�ޤ���xŦ��Un$e?���in���K� L���Xb��K�^�� b�d��R�%�� Y�S�1��Ա�&A�l8nӁ�-��tͱT�dj=f��X�ٜ&��ֆ��;����XxNB�+rɻHo �Rw
�\��4�3�;�}����j���81ΪM�W��E��C�6>�k�4�'.cttP��s��+��|R�)�y)��rע��r��g�����Z���}yy��r����i�*� �Bb�
�%qn�S�,��O�6j��L%8��6��?�Sn�8�?��9�p�����WdaJ�^�ۘJ(�:�F� o�#@��wG⿁2.�YTA�X�`T�	d�g=�p?H�7R�ŭr���.,��}�������%3%��鎥� [�X\'ZI$7���y�DS�	r��Q���$,ʎ/�c	i���4����BRB7���Q�c�����Z��W��%��R�S��KE\�a���O,��r����I1P' ���,tT����|��
�$<�؂��'R߉_�+,�w9���bɖ��j��Dن8��<v��e���	0�ٹ�I�̓�U�QO�Bȇ�Jȭ���Uj6j�z$0�A��Y��~��X��A���AB.� >7U-���U���h�U�j@�y��W��^��G�)�#�])涝��f�E3*B�wzNq(�E��>p?a�w�k�J�aM�	��`3'b��!�C���}L�\�F�@�9�;�����S��Ս%�ߵ���P��� �JE����f�V?eۇ�W� ��vF�soɃO�H�֯0�m��A�yֈ�i��k�Օ���w�����rf#]�@��CL��m�EOӣ%�:��N��؎�9���沃M��V>d�H1yD��&��E<���3U�����ס�ե��+6�=��+����{�r�QZ�ބ��sOt�f��ȍD(��@��{���j���j���������a)_�fo��ڡ<SV}����W"� -�
�\��ڶޖ��J��}>}��q8�gD�n��5�T�(LIu�j�����㛷��it�
\�o��C�ˎ���o4-�d󂬀�
�����Go�`�J�,��2²���j�`q��ɅU��~e����g|m��\G1� �%�̨7���4z$E�
�VI�zs6JE9rrT��ᐦҰ�{��+�xپ�Yʙ}��|�D�[6�:)p�(�4��8�|�}�&�4�f�J���2+6?���x�	���e��c�4'����)�9����w5�xi~'�+B�W�mFZbn�3��HU܅��2� �Yb�'o�[�W:���1����9ʡ���՛��#�A&���*��Yy�p�΋�qR��qG֢�&�Q~j���lW�ir��w�f�ﰏec+9^�7�RO����"��V�.����L�Ά�������\���hN�P��
z�S㕼JC�o��U����0o�ߐ^m�$���Ǭ�W�F��͑G-n}�̜��\9q���,�R�=.�������vv�Ƚ�`��ncr`bn�~���k���1-ɷϭZFc�3���1����zud&6[��͵7i��8�����	����)�`�j�Jik�-�{5�ޜm#�9_�B!�L'�W�)�O'̃��- �}~!��XO��f#�k��l �l� SC�~Њ�me�E,��OI�u�i� ��jN�I���b2n�9~�=<ķZ5��f��N����	x�2�loJ������Ðv �N��}s3h���/}��?(�6�[0�m�+�Q��|�B�&	d����~Eـ�浛F�15�~:�>��p,�f��W�%z���⳷hd�`	�*��}|mC�?��	���l�5��6���ɤު��V��}g�Tɣqh3#~<"-۝]�蜮�۬sk��=�S�Mb�r?`��Kr<$	1�B�^ª|�P�������9I/;oLώ���˒�u�^���H�E;�������F����JK�*�:���ꚽ��#%�����T��s�v�|4]Q5���������͂�M�5��5]�y�
z^DA��pݯ	��ر�_k0�,V�խ ����F9~5M\�ឳP�"���@���?�~�ϗ{?�">+'�)��~���q�w���.�~b�����Doj�)Ġ�W����
�K�T������Y�"n'�T��b�/�=o��W$yN� 8��.�&�x���t��b�ȟ�ی�h���>bדe�'ޅZ`6y�#�y��1]���JuR��B'�4��kP��!�� �=D݇�}v;�
_�ɕPL)�W����X�y\�S�x~�\�ʮ���m��[��G��\��zg�_�,�/���)�����[��D��^�Z]hc�-��,D'Gal�@�5I�,`���\�*m��8/
���w�:�����SW[l�����R��@��N��x�?+c����d�a��}AZ䓭��|�*�7HPAML���R�.�!~����kYA��MW�)�WG�L�����ʒ��K�Xdt�<�a��4^I��\����&\#��`,�\~ �V�Β��yB�u���y�;*���I�jM�� \��%g묆&�<��(H�/[6<A��l�dU��yb,v�b9�G�������^�Z�Z�X�����r��sY4�k�ZC�x�� ���Q���*�Ư�oBQ9�i;�gByyH�$0�P Q"�/��~ˉ�G�'Ob8�7&���b�֩Ν�L>�M�^t�2�Qg�z��%�a��/��$ۏB�'Tp�H�������k<<�ʳBx�� �Ɵ��O�WA�/X�1��O�����i��|o�R��ދ���� ^�bJ����J͝l���%۠P� �����Щ{ǌn�,��a�sK涝I%jr��l�Ӳ+Us�Z`�q�yl�3��Cv�@��mpn��Ok+Vy���v!�Xo
@Q�Ì\S�&�ϸ��QօD���=��c�=
���O�0U���s� I:�������7����	!�EƜz�2�v�R���	��I�Պ���C��'T��&T��_�ifS�Ұ��jO�V棧+b� mfloC� ᧶[u����7M�M̝ul�w��J��i���=������ȯj��[�ըٳ�h���c�b�5zZ�Td���f��O\�? �)]��l�|�XU����A�V��>R7�( ��R|7�D��Ӄ�5?
,J�e[�ue��O�8TPl,^r �z��>����45�����+>JI��t�����*(� �~wt��ǽ��ka �fg�f�~tȤ3�J6��$-z�e�K�B�cU���b`Ɍ���~�MC����b<��o�}��a ���Y?���ɿ�1+�����[� ��^iK�;+��y��g���}c��q���<�*т�����n�{�W�Ix��m�H���Qj�\�-a�&A6#�ҀqPAnb�3�&h�ۢ������je�lvk�@��_I�y>���vӘ�R��d�,��p|[��s������[�硆�j��j�Sq�*�Z;׶�c's��	X����.*����Ta�>ό�s���ԫ��N�����5���T�5��e�y���^8���;���+��V}DJ4�c��P��W
nyr��� �v��Rn�Nz�٘�:�����d~�� �V��R��𒮄&^;{\�[3<Ǧ����O��-��b�W�6����G��N�bvӡ@$���b^�/�L��A��]wK�x�P+�ڛ���7䑺^�wY��}q J�J���k���r��S�>}>�[��dz{΅N�z��|��Âȥ=��	�9�}"谔��3�L�n�Ģ�G�K�^��f٥�}�դ����+�YB���Y)�F��/Nq�:����Cj�.i�>
X�#z�,9��&��x%�L,��0\�DSX�.U�R�M�X� !�����!P�6��Qg�/��U� ��"n%�6��̩�j��?9L�g�~c����Hb ޝ ����ʩ�g��
�Z�^�,qӋB@�V�N�����rУ��� @Ɍf�k����.��I��rPq�W%Z?>
Ҩ��4������s9�e��X{#��+��j�h��'�����t�-���nG�#�K�;�e" �O{�`�2��P�x5���pʲ����^��F�n�Dwh���W��W,*��W=����WL�g,U��j2�1ᰜ�@hӛ n�6l�Xr W����K� �];���z��W���}t����9-�<V+o�����E>������� h%`AV��Ű�S5���i�4r��UT�����\� �y�E�%9Z<`1@��|��r�&�T+QdQǌ.�]� ���"��<i
2Q���i�y�7����O�h��D/^���S��x��`T��w�vg��$�R4�`���X�)��Sy�!VgЩU�^D�
M	�%������[	hT���@��
����܌�W6H֡2&z *?_�-ϷB�7���? ��J7g[N3��n~��GIfhrԹ۷0��U�p���˛���<s����򱀦���t<��@����NCK�^+�I
�~jl��@Yǉ�DI��"+7��~ǝc��0�,�-�I��`mh��H~���'��X�O}�yTI'���[A�=�`[
��H�gB� _�s*�&�Z�!-iP�%�֐�]Jg��ܞ	D؞���F�M-�?WwxS���z��@��a5�D��]D������-T�&����:|=Hie����3m"���=��ƕFM1YK��[Q��E	�Z���*�fK�&(�%���u=)eieB�пZ��ђB
����z؞�A:e���9���8�s����I�� ˇ�|Aсl�yB�(R�ԋ�*���gr�5%È6$W�݆j}f�8@ւ��J}������O��K�Q(�'���,��^Q7��,
W6P[��<��~o쵼��κ���NZ�7�x�ra\ҷ'q�r�N�Z~�U8�i( ��[r���Rq]��8m}`	h  G��M����[��-�M��&��S���0f5hRи��l=:+k�-���FB��R6��_2�洖CXG�-0D�^[m�`��#?�<��!?X��J��6���ӂ��)����T<F�wX�+�>�eC��zꃹe��=���RZ��*tZ��s��	l����r?Bj�+���C�6Y`�Co�8N�y���y_�eP$��bv��I�1L���e���=��[3�޶moCc�v��`��+8ɛ�_/����5�Nb ��6�Si��<���C)������*F^��H�`g��o��@z���%��Kbղ1�w�>)}Ҧ2I/��/v���=��	�D�o��P9�&���j�+��,~e#}����&-��u�&�xP������*�j,�������ZD,d&���7$W�r�N�|�|UѡM2]`Y�,�Ğy�a�-Q��Ju������*f����J��r�S��"=��UuĽ�����/���As;٢.�	��J0�,U�^V�h.Y�?���k0�{�jQ�<3�(�&���$�.V�WD�{abh�3N�v�6L�Y�?k$k�\oQ\7T��c��_t��׈�E���%��8>���`�fr�B`��%P=
�3��[wI��Kw��4�*�`�(�09H����g��r��u�@����JI��
/�.6�=�)t`i�nW�)��J��(2l�\PC1�c��.�!�����X��$�;��=8� ���3��v��cv��sh�A�,��z�$����d���}p���0l�g.HI�a�X�Y����o�� ��9}~�~������7�td3+`F�':��@�g�1Fz�����5�'[%����tÜ��d�眧mzW89Aj���B�Z�������g��%'��\�u�m�2��Na�8�m
6����}u���Q���τՓE.��p8a�4������dg+�׀$�;n�U���y^8��U���qf�ލ3e��Pe�0�;W�tyjD�>�rku���v�b[G�:O}f̴ ˟�B�����{�NPs$iϮr
L&;��]�2X{-�^�0����x�@�+�sܨQ�������
�T�cfr�U���g�*>��E�%xdfk��x��qj���󂦻a�5X�`�bZ���9��X-뛇l1�8^�����eux�"��g�z9\v3�  ���T�j�E��_�ͺ@�+dڸ���JxH�GA�N>^}��f�-Qy[�ShϛL�ibbo�oF�1\�� a��ݲ��z'�t��ܐqq�Oҳk��d�dǟ�<�ka� w\[��DG��T|򌬏+�5��窗 �
^���͆�V/���~E�D�TF_�-�:"��{[�Ʋ���#5Y���� �M�A��@&���6^���nsxЂ���&��I�bp"��a��:N�T�=�]ɑ8�e<�⼯�2k�����d�3�ݣ��]�|�ɌM=�ܾ[�!�[�!_�����Y)60:6�����w���z/IU����i/��@u�c�鶔�jY5z;�Jjο$0oB�[��`.
E�I�\�]Úk�|h
�ӣ�<΢��iA����sϷ^��J}�Cp&\݆>��Υ˫Ӽ�։+99Fi��~i�����D�G�`E*Op�:
�����KC.�eDc�\��tݕ?�zH����v�T:H���͙�(����ncy�M��7��s�q��<��1YB�Xz9N
�ژ������j'�HwJ+�!:�p�zm��:��OH�84����6�E2Q�t��MH�RҠ�e�<Z]v�%���+"�>p|��F���G�*�>4�1���8��_�ɥOT�Ms�F�:����j���)D�B�G��_E�\*�����1+�C�:��Q�-�K/�O�ͅ]q�.$sn�V|�봣l��n��_t��u��ȋH��h�3�N�&ۘI�	'i%^?��\#M��]�w�H	d~��l�����ޫ��U���Gw���ɿ��Wmح�\GʚK����&�����$��"��0+c��I&�˟Y�vt�:3���"ߘG�r��U����[���ח��p�����Pc= #zٚ���G��4��HS��(y��9sޭ�`���d9����m�F���Y\<����	�G�X�7���G�h���c<��S�q:z�I���1�'De�c-B�I'���5��K���^�3%��-�	�
Lɓ�MH�9&=�6b:��Ӯ�ST�EFl�Q���<@سSl��޲�?%(��~�}��F7L_3>�5�u���4}�<���9����e������
��-�XUI�b������W;R��Ȇ$Zk��<�*&�Q�t����{��韡�
AF'd�=h��D�a�`a+�`�J8'�a�&m����]�����*i'�G$�#���0�5�z�����y�"�J;�;���1xʕ<�a��5(�p�}t'_0��Y('�Tj������n�b�ؽ/�ӧ�~>��G���?��w���g��}<��݂�m.�	w�$�5q��EDЗ-+�~G��O"����z鑯���m��ix���ֽ/l]�5�[�h�{���{�����ƃB�%x^�!h�^�z��4�����[����D6�����,���������]p�I��}�X|ST^��>'tR ��b�?c�KV�T�fhɓ�_�z6����-��i���DD�^���8_`;��;�RF����Ȉ��D�j�U�vg���&����u�N�AVxR��V�1���C�����P?>z���5����_ ��N��vu� -�ޞˌB]�E���֢��*K����0>���U7�i�٤�V�⃛�"y0��ب��� w���̷�ɷ��S�)m������T��G�g�/E5���F#�������v�%>p�(H���H��s2�@�O,���C�^�$�.1:�����J��l���
 ���Y�;�3F9�%L�y�T�;��^,�>��S��a�W
�U��4��ҋ,k�1���DOՖp��tq,P����H[|�v�VC��_=ّW�����vb���������T�t�!�1���kDW�/���cJ^JU�/T�>e�9��O1�q���E����(4�p1���j��!`u�4C�*NtY�C�A����7������(�א�pB��A?R̊��ٍ�u�S���H�ߎ�}60*W9��A �32c}U+�^�9��D�J
�wF��(7?C-�z���
� �1o�,�ڤ+G���m������)0��f�S�)�@�;R���Nҕ�7�r���O����oir��F5��*�Q֗����|�7I�1|Lf��������;÷�S��{��B�T�+�Z�m����7iF��.��%����8 c����u�0�ZV��HgO\q�g�P��ѼRϘ~-�)�}��=Y��.�q�)kk�>�������J@��HS����A�O�� 8�'w��v������0�Ĥ$�$��!���Q�l����b*���Й�Z*���������� ��x�d'�޳E-1���W�_d��������%�o��&}΁O
��_(d��D���P��@=��C�ӃMX
���@����#:V�&dLa
e�S� γ0�y��r�K�����l٦�9AC	)1�Rud�;�H�t����ء�r4�Ą��M�(�wk�&C� ��I�B(a��7�&vR�Je��ff�g��V�ȷjh}0r��3���Ug�äF��Gc^�|%D�e�n��@(����)����O����%� 9 ��>Y���{)�4"�@5ǝZ������{i��$�����g1Lh�?EU��1���o���?���i�� ��Q�j4�@R����\����@.��v�!`Xf��R�b4Ƞ�j�sk������w�ʚ~h@��,k*Z��>�-�� 4�.tB'S�[���1������A���),]T��f<���{Z���t�!|n�R��O���#B-�g���	�r��õ��Rدsq�]�p�j��	��Jf�su~�m��N������Z�ڑ�C%��
����fV
�R�С,�w�j�t4�`�G��BKU�]�שV3���^1�Վ�'趘���%�}B��y�:�ʰ���<��C�-w4��U���"ЇA���sw�j��S*�6������o������?ŋG����&��B�.@�Rj�_��Q��	���:��yV{�O�,��g��\��e�����
ӗ$N�<#+a��"�O8A�U�_��Q���2;�r+Li�_3�oD+�X�S��h���0�X�fp���C�8r��v׻~�G�G�*�UB�׸d豨t ��r��e�AeTZ�����^a�i��]k���Q�ޓ�L���
���&.ookz@�d���khy��D�_0�@,Hf��$��4�����W}d[��"��o�?֧ ��#����8��i[Tr�Ӽ�d:��-��"�g����R�+���,�H+��XL�����ΜD:��-���H�M��&Mu��/�o5�?��E2M�(oy���k����)���/�$�
=�d]Y�����k����+�'���(d�XiK�G�} �H�Kr��wzɒ5�GtѤN����"�T9[hRʊ��ИE��P� ̵�T8�(���	��×��p8#}YP����1���� l_>ٛVi�^}k��+6R����zX?~/o�Q��P��k�_:��1��5t���C��;��kB��L߉�唸�	�q�.+�]h���V����s�}������=�f��3,�� t%���^�_:v"j�����jK�j��G�R�Z�+�T]>�J�9��*�Fn�m���ν&@��� Ɗ�g��AOz�F
Ē@3��A�8s����Fn�O��#+E�(�ײ(]�u�T��[���5�w�}7nEm�ңF�C0�i���#ש�c#�e���w���=%�רJ�T���K��!��)�H��B'!Og��4ӱ.����&�"R
^�8�dRO���TNyģk�S'����S���3���
��
I�(��.0Q*F�4���h�D98!�
�C�I:�T1n<l�V����H.�أp�6�����������Y��W8�ź�ɻ�U�VELѸxU��3=�Dn�x�bH�Ƴ�I�b|�E�1��ѣ�G�R"��p�b��k)6gC��+5a���O#�w���gY�\N��щw�����A�E�����F�pX���Ir����i���*=�O8����T"�.
�wR÷15ҟg��M���1�Ue>c��(�b�b>F��m�#Fk7��z�"�)cz�H�����u���#C��|þ=�F_�r�I4j���B�n2��3�&��<�7�U��P��jSu��q�2�{y"Г��O�����XrJ�>(`�o�@��i`�)#���(L������t!��ݫ�Ɖ�G��������ܬ;` dO]�aPW� ��]!i�L6��MK���I��䁸�7_д�%�i�N14�7R�S���g��~�xg���5yc
z�cP-� ���3ݢ� �l�8@��w�A_ͬh��զ��/��rU+����i����@q�"��cJ���;�+}�v�
�0��F�3��F�/t�r��섦�/rfگ�� *�C��	�,&��Xݦ�A}-%ˠW����Y�(�o!O�Ʊ�?�j���̨�o!LP�}r�7Ոn(���a9dw��{�(�@6������ϱ��c�)����ev&գ̻����ϖS?�D�+���C��]�����_$xɠ��)a����'��>��*�(��g�.���䑰yzT�z��Yba�SxI��q���p�抴
�dh��W��k��!ї���?ш3���+��?殃 u� ��-�"-@�p!����i.��~�a���]��ͼ+y��rb�[��c��c��a��I�C˜��~&U�1A��L�3�+�k
� ;�ߛ��c�y�H�&4/����S�}�+��NGx֝�3H�Z8}&�2����+#}�.)�4/рᓡg�<S<�=Ϣ�O����4|W�J�	Ӂ��J�Y�g��F�^��Ŋ���;<�>��ĀɹX�z���8����>����?<!���]<fL�K}#�)S�wlL��CC}Zͨz���J����%R����S�QwW���K�VX�($��$���,�����{ �{��/m��Mܱb^���=
����G�Z[/��]X���9$ɾ˙��Az�[;skj��"6|ɫ��M^��c;�o�<���C��<#H���o� ��������co*���n���h�۬(q]O��d 9��.gS�1n��#m��)��k.������˶p����(Z�*a���c����/�[ʋ,���\D��޼�E�DҌv��x��=m@��P�Q-� `��u�۰�3�n��A�����kT�X�,%�C����(���m17pE���?ᴛ��̒O�����1l�޲�^2%��zIJ���c�J�K0ο=��`o�/ܚW��IRB�����X���J�ި�jn=	��f�l��!,��]�Q���p�@���!���	Ue�/
V�ҐhF��i��)a5G�D=6��bt�w��U��L(Y�^�
�#�V/ȫ�Ԝ,�lN��cJ�����Mq޶6�9J� 
au9���u� ��N�Vߵ#l�a�D��4q�Գ��t5�*��]T��&�qȴ2�|Ii���q.�\~Om�	��i[W&\�3��r�'zK�����86�pId�J��Z	��<�������BBUYF&.�m�����3Z�K�vrq�@�r)�-{(3I�3����
$��#��g ý���Oշ��\l`���~�z�LY�)IE8�mY���5nct��R�Dχ��ɗe���,�^�V|9Ԥ�1&�?����1A�簵u+�E
W��=Dzu��uv?>1eP�/2E��˼-�t	����<2�:]��)=��)[V��iu��IE{�h�J�Ƴ�K�2*B^��W�C���ޅ�qF��N�eeF�~j�B o���D� GL�����
U����ıSbf���|s�x#��r��%��^�
��i���>s����y~�*kݚ9��c��.3�,��+ߠw�Y��G���h�0�C�9�*f��0�W�=f�\6���ի��&,�ڨN RϤSd���e-љ���An1�={�Ł->a^���!�Y��jd�7 ��fv����GV=�E��f-��N4�G����y(v�'w�)�of�S0O�d>���o7/Ny#�q��1%�H�Ҷ`�C���M)ޔ�@�)<�J {����T��1�Y3����_!��U�r�S�f{a�θ�Z�u1���G�#����۸t$��)��I/E��\�d�&a�8��e�U;eܓ|Τ׳�g��\��"��	]�`���^�U5�a8��5-]>��?��t�$u�n�b#��5�[V��>ª�X1���	�u��Jw4&��b:�k�t��V��T�1Ϸ�+�h�犀�c������9�j��ґm@Izbw*o��@a���?@I:6H�r�գcL�下Mp�
��k;G��"C�d�A��v*��l䒍�n�F+ {�9�'�%�@��J���2˟|׿�q���v��~�^m��)�䨲3�϶
d�凜�}��i�d�!�˛�H/�3����_���?BČ��=�>ʧ�pك�����2F���S��CC�h����g�� Q�f��j�����Il���LώT$��b�K�I��tZ�����°��Z��_Ԃ�R�|I�M*��`�M,�CA�*���Y�NɄ��?��8-�2[����z�M�y�_ ����-5��3N�qy�쾟���>��j��~���@�yC�o>�Ǣ�`�F.&^��?�h�Ӕ���6rK�>\���G@��;a��~��X��MxmC� OroD��{Ok��韠�93��9�ɲ=��P���Bf�'Ȩ*��<7����Q�\��~�\����́�=�Q6���ɐ��-kg�1
$Ѱ�X��wJBm꒣�_	L��X��G���dP����k��t�D
�dB�x�ŗne���3RP�ӌ�j����r9�G��ۡ��߬�-��؞`��}�]!©���=d�կI� ]�Ďǜ�"K,���
ɼ�ݼ<�Dl�Z�����[�U#�����#��+��v<�r�۬���R�����̂:�������AR���ba�u6禊����͊6 ����!��f�z�']#��P��*�ĮW!��\Mi	ϩ��0���YQ��ӽ��}�����	��M�>o&(��w�m=��&E��+Ņ���{ؠB7�]Y>֜�~�?˘\��s�$�@���t6����}������x8. s�VN��������8�������;b�0L�	��hv�|�ک�����ї�,��ܟ1�^�F��Z׋3�o����ٹ���U�!�a�����=��͍jO�_�mL�fV�d��/`�Q�3�A�9��C�-�N�� Ro�
1�ٸ�d�P�W�կ쵫,���+�f(�1j�Wl4����cO�����_?_��{��0��IWV��c(�yJ:͘��H0�N��Aoewl��¡^`B�j��!����`G�o�!c�������Cy���HC/���N�w[�s 1 &�`��g$׹c�dfڨ��f�z�IP&����\z�Þl�4��5��i�%!��o9L�j\���ߞ4�:�F6z;�M�Y�������Q��5�QJ��Q��曰|m>8O���go�.8͐�`�W`�ɺ]�)�9�Z���m��Xw�#l�9�wӃ�����K.v[�+,�E���#���P`[źf�~_�B�(X�W\���B��q�L���#-�p�3������h������Q����� ~*|�pK����.'�1���C�)�������4��<���Dbz�j,�^�$�%�Ul��	�϶Z�!�+S�|����������*쯎|`ٹ=ٞ�blĆ0�$�e��YS|�o��E���L���)IR<�Zࡶgx��4���G]�����'��Gw�1Ce����^��h�R�SA�,>��G߱s�"ڵĪ~C7�&���4�?����,��bf�d��Qưe��p��+��:�z:�i�Y��m����ϼ����J��g�UX�A�`����f�M�)x�~t��"�nj�1?�O2�=�� a��z}���9�3E�ػm�_��a�����Rs2S�٧���,��OrV�Jh����U�k6�&0�0�xO�����X��r2�9\?���L���Pk����d�.�k��ׄ�p]®� ���A��kG)���4�������@S�q}��3� /����e�	��^���X�0�4�d��IA���6��<�(����c�Q�u��T� �Y���-缦ޥr<��g�!�f��<J�
�����*���P�s Q(�K����s6�+� ��}z���V���=��l~D��mQ��U������^�s�J��\HNL�Ҟ@�*S%M�<3,Ow4n����,s6�L�R\�GiK��k�C����@�u	K-���G�J#+N�W���,翰���I���J}p��-�
<t=1����	�J�&��r��i��sZ8Thg�%�W���2�C���A���|\6�t҃R���X�宸�|i7B���c�����V�8q*u��dw��w�1�l�����9�[�xC�ϊl�Eyߜ����eD_n���E�UEZ�^/�d��#%⪣!ǟ���+71��H&4幏�׎f��_��ጼ���s�]��#�&�Z�S;jm��@(i^F�*�S������{�>�r��qH�c$���L�}{�bֻ�yN�����p��T��g>��Ԙ.��H�\�p^e$�9�ن>?�]r������9Z�Q�V���'OZj���/�/����}���<���J��`�ST����6����r��^���#��M��*p��h�
z�	+B�lJ��"@v�ʞ$��b�̒�߭C�t����B�Ȃ&��6WR!hd���!��Be]�-*_�z:{Ծ���d��]���މ�v,5�0�����-�*�������c��3�uʂ���Yϥ�Z��Q5��?M�	!�z���`�!ڈ�w�7\:��7$��&��[�W� i�>���?�7���Y�0�����s^K�+�Ʒ�`Y_�����*���kDo�R�a��\�JFŭ��x���F#V�+����>TJ�[����H�>*�3#e_���?~`}r��kC�ך�	 �~4�J��6�����%�(���H0)o���YA����+낆Ώ���Q�q�V�^��O���yC�*F�b��?G���h�a��U�"����>�]�����n����i�;KxK�#p����#�B�N,	�b0N֚�m�f蔙�g?=��^\�Uo��\^��0VU�ˆH;��#Bjn�a4l�'e��d?Kٮ����R��/��nP״N'�?aa�8۴���B����L��n�+���F7�:����w��W�KS�o��c�fԖ�Ӏ���1�L+&�w=�e�.d�v%u��k������nk{�!��U�f����yw2�~o��2/�-�+�\6�@����	�MuT$���T����8f�B�ӞN`O���n��?Y�<ck�B����!<��kրѢ����|H���q��n�%DBd�G�Q
,8����#zW[�Dsrݩ��;�CBfap9�����ѰN�����>F2��_��(��6��,#�^�m"�'��|�����]0 p�=}>����&qh��Tzd�S�o')&Z�߮��_�й;s�2�k�5�#��?�<�C	A;��oT�b�эNd�g ��ȩ.�>�m����!�LW>�Ji�/�6N���q>����V)����y}P���e�y)�Dͺ�Q��.@��gw��$!���T���Tg�&R��s/�ࣥ����8���TWġ�����Z���)���\\vk-���2��uv��[�|d�$07{\� ō9<IK�.4I��>���S� �i'K�+D-�<��:���ĭC��H[o"9b'Bv6���D#ʁmH���~�
��@wgI|�ժ:���e����P�"I�%�]�d�$}#pm��fnO��b�����hky��r�o@���](h�>���b�;��=�C*Y���ԣ}�V'b�� �!�T���$5(B�������jk�8�f��OW�����6�A�+`g�԰�3�ֵg��8Q�,��Ψ�}�o�q=^v3f�Qɼ����:�*|���Џs�AV��P=ssWD�l4����{Tf� j�7^Dt�
���&<��G(>6��?>
�lV���E�-�5��Z�>!?���h`��W�;u��%K�z���"�v)�U6���P�\�zUi��v�xV[��Ҳ�S��Υ;B����l?Rz��Ϻ�{3L�xL#�m�h	�)���2>4���(%��kR]0jnش»PU�s�*�Ҩg�I?M�T����ѻ0a���~�/���!Cӊ�}c���E���`����tH��K�vK���;�n��92�������	}fJ:��i��p�<]�.���0�f<�pB̛6�>IOi��!���@��F�sͱ
�5R����sA�t�� )�ހ�ж��|t��J4�ܜ�H��!ci� �$��WOĢ`�Op�P���M�0���  ������&����I��x�t3��t��~������.�U��)h>(����w�<0A���:������qZ���HvIe�	����*Hm�ĸ��!�9�