��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+�������;���ȹ�v{2� ۝ߎ#�W�ӂ����ݠ��>_g5���t͉□K2���Ec�ſ��`\_��cW��Y���NB��*�!�#-/�����0�����e	�.ZDG����g/G�lз������s�VS�]��	�_,��ܳЅ2꩙Ō��M=룯+�&HfUk�@��%��.���cm���pZ�^�&]C��l�QQ���UicM���*�qz��ZU�^u]�2�=>���J��מ�#�^Ķ���l�\*l^���F��A��N�QI�������T�xĞ��pǚ z���4��)�7�z�wcl9du�f,u���� OK���ي�H�I� ��l��.O � F�		�,& �����ͽ�`� 7�(������,\��S�!�4��ݮW���l@����1`q�f�>�U�g��E�����a�md������N���+���+���}���t�
I��-�&���I;c�C&�Q�J���5땕�?�Z|D�YP��e�|*���#܉B,��S�(����L���͙�p�&d�d�d;B�Hᨷ�ǻ��qa�+���  YEɃ��)=��������Hr߈�/G�S�>������`0&	�wu^+�#C)H�C��f�k��U�lv��v��״KOgC�Ѯx��X���8�xh��]�
�J\:�68i���Z�O	G���[s�B:�E�6M�x=	��Y�hw�946�֊0�緪&�td����q��)6�wqx��L53e�ș@h)�}Z
{�z;�L� �HW�o��>�������T��Ք�x���W��#�϶�s��B�t~��%B8��S�96C�/T��C<����!���:o��T�v�3R0`j�>��V阜��[���EU��J����dL/t��k,`��:RJ�B�I���'�9)�@j3VӘ��Jzxf���:�)��9sJ]
cm �04�S^�"�_u�չH�]�����<fYV�.m0_���'��č<����'
�pCF(��c 9�D�6�����7�m~e�����lB+���^A�΅�ǫn6YB��\Υ�+9��//lz�jp,C��~ވ83M
t;��6��\m��v{5[3);� i��
"b�x�᯵�r�dj��\�#��t��Cg�O��:��1d�m;ԟ2Bu��+�c8���ҽ�F@�؀4�@�Q��qW��.'O?�y��x3,;���/�� ����3���4�����Q�̋�CA:Yw�_v���7l��3���BV�� �@��_�5�I�YMPh�rFh���^]�+�J���U��Pyq���,yЬ�f� D�+6�e@�*�Fm��P�����Ͳr$���b�?C�1�X�͜���-�;Dt�@�)ff���@�y�h͗!����u՞* ͍��z�
b��bC\���V�o_�{a��#w�6B��}$NK>�4�Y	|.�!�_�%3�մ�G���:��ȷ*�C��1/q/��}���^MXD5o�hֆ!%��z��EY��2�(�:�±[(@��Q-��t����Ҟx�S`#[�0D9Ewȝ`��-�Z�����e�=����xL7�=̦��D
�S;�� �cF�m�d ;J�G9a��B*Y��s���>���%�'7&����!�9�f����O�2���ޝ�0�ҡƗ|,ĕ@d6��
����ʧ�@
�e����t9"�c"�?i6:�1�P��4�ԯ��������V~���Ķ9"V)�*�/�^�M-�r�����:�*���[�ͩ�;�|�#��J~ �y�-}���f� �c�V�Ed�<�4Vm*^�����e�x���e|ﰱ����G�����dάVk�ՉnT(���V�I��WͨJ�-e��wϽ���U��GBJ��ň,'�n 5��?�An��L�B&ʪ� �m0VB�y1"&FL�x}��u�(�?��aK��χԋ�X9ߺI��~Z�ս��ڭ�ma�%5�~�X#)��ݬ��eQ��b�"o�sX"�C~�m̚�3_[�O��2�G� �o�#k���m�m��w���gf�����QE�~򃍀v����'6���߮Ez]3y������l�-�����l��c���Bo"���.&�Uuq=�;�{��rTc���`	�Op�V�`��f�?�Yb�V�u?P�����O���J%�3��؅;�Z�B���P}��$<��)����4ц�7\�/��Z��<s�j+d�\�i+;��&N� n���t�O|j��`X|�b����C�4�a���Ae�P˶I��di�XD�&��/z�ynϽ�{���d��1ǳ9�x.��g��3�͹���jS�B����GC�yCy���7z0��v�%�̘DKkIeI��4I
�����k��uF�hq�'#������tc��O��)۩�c*T������b(��X��%Uɺ����k�ꘖ"��-���F�v1ow�T�|�a}Pn�JXa噜E2�zMn8���ß��L�������e�m�<��� ���K���d[c
m<ܖ �h��x�h����~�[J�bP^�p���$P�&P����m&t ��,y�����*��?k/�ԂS�a]	�.&kE�k��2�zyi�i En>q�p��H����'+M�B�*����g��'#L��|=���+�}T�T&{T��VQ�<O:X���L|�w8mv����$K��t�P}�S5���F =���ѸF�a���y��:�����<G���hfg,��}|������տ$�D����.(E�_�Q�I��+~�QX�K}��2ZZ���I.`�_�"�4�Ϯ�W� b1�Q�k�~��OJ����� ���H���i��LU�����$��n�`�E� @�ۑ�$QKVV�wn���r8�e�~Z�Xؕ!D��@�ob
B%�=�
m􄦃HN�gQw۽�)�jZ�$�a���X��T��+(�j}�_L�Qa?��U�Ë���?��®�����J������3X~~B�����Ζ3�f6rR�7��~�n�I���G�Ҡ[�	i��&���]4(��ca�e�)&��0��J�KlHld��Px�E��@w���P������@:5���7���\�dúK��h���D����ym�iωD�{�J�G1���� {o'+ټ*��~�	�*��@V���D���yM���M6��k��[�bD����7�I�{��|��B|�%�=����(!R�v��*���.��P�]Aj３��l� T{���}܇��d+g���v������f+�� ��m����p�$����T�i