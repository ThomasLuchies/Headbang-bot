��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k����W�z�N��VXi^�p���d����So����SaL�X�ģZnHt��ҩ<���@ȸV��k��Y:	�|��.�<,�'�ޡl�	��E��V�mo�_ ��9�� UE�9Ĩ��T�w~�uX�i<#l�Gq@�D�6';+���U���W��0"�FW�D$7@5 �1��ݨ=XFN�r���T.�NWW��^JzS�zğ�H�`[�Ƈi���-��xF`a��
�y�H·}M���`m7�M���}a��vll������.�.G���_�	����e�����꒲��Q�!� �Tt��S�P$rұ��#���
�	�"��^W�Z�0����,����� ��U�v�Ϙ����F(J�z`�1���H!*�a3dQ�?��iW���I���,���{<qƨ���X�t��sj��a��?b�٧g�v.�K?���	�w�_r�x��B��t��I�����4�<M�������a�{g�S0��U�̬�7�j�!*���3�C�OB�Q/���K!y��iX�s׿Дu��C6|9}�����=Mbm����K���>.�c a�݅�8@"����F�N0^[��t���k����#l +�>���q�x�5[s��Ǘ��%�9A���,d����j�
��!b�B�(�?:\'����;�OuMe��(���ϙ�gZ����QO�A�H���&��8��w��E�c�Y����j��dq7�@|������޹��;�	% Ҟ-$�=��gvU��'B��0Z�|H�3+H�2{�ˌ��F�"��֦���� 76��l6����Q�٤'�_��c����O�t�V�y��������$��T����������-Nkʋ+/�X�e��  ������[$��{���ó�%בW�H���B�G�������BJ�? ��H�)��SD����0=�)�3�V���C�K}�4��Ql�,C�m���1��������V�h�In>���QHʆJ�ݛ����}צU�	����M2_Z̧c���Gy0�����}s~hic�ٸ��󐜉��pD&�����}����+[t�'r�0ո
���>1�ڽ�Ό�{.}Q������<�#�� p@P�|�E�f2�w$��d��|����UQ��RK8Y�{(����Q�$s]
�M�˓�KM�Z!#T�3R��@�A���s�n;b3|?zi�	���U/���֕~��щ��������6o��O�uX_��M��
��L섇�ȜZ(͍�,i���$e�sn�*�-B��́7�N�o��.����"j�Iza�N�R5�*�����!A\b������a��w��S}r����yw�m��)b�1ܼ]E�w��V�����a�Ԫ܋�%��]۴���M
���X��+�	������
����ڂ���c��/�4�G��S�x�L�ț����Z�&E�Z�2 �u��B=���n�o���l��=�eY��C�y�F�=7;"I�8��+N=ʽ{�&CޢOpW�ہ%�r�z۹J�.7V*�@�uG������W�v�5��5D�K��6!qۄ�JvPɤ�I��cݩ��˰�S����⮑�s�����L���=��ٯ|�d�� ���o�|�8�ͳ�P�$r�پq;��w3�T���꛼w���J����"���줶����N�}=On����4����D���Ӥ�u�+WS M����@BZ��[lew�DE�c_�;W���x�`�r��EЍ��(���	�׈�!�5���~r�Y����\��pc&� )�{D�K&\3*�W��4�����-Z1��p	���ݟ�b8I�Xw����߫�'�_�(>��j��X����SaSsHaxs���],��-fBMH���G$���b���ڻxg�>�GԛX �&0j~!�Z�:E����"/A��LE`Ic�h��IД�)�V�j��i6�t}�g@�-3r��@ Q�/%��W*p?']�X��Zc�w���D��垭��6JT� �_&	_;n�'����y��<7�1�(� ;�7t'�j���ú@G�:����|�AG��S�ǡ����[���{f�C�� ��M���V � ���M�8 R����fr�:'���j��}����A6, �W���#��"�;��@W�P�����Xh)�YO�0KQ��A*h�N���8�-W+
:}�9Y�
�a1G��<`U�9^�oǜ�"n��8�	{�����S��7�PW�j����X�.ia[�2�0"#���"@�o�5�{2�s�q�C�E�[R�zk�C,v�.a��AI�Z͈�2�s�u�d������y��7!�-�!�u�z���/b��c)��Ѿɝrr#<곬�sQ(�?a��=KYl*W�I˯`�i ���wh�����,�G;o�;�ф{	�Pi�9'K�>I�S�����^�����VI-}���L�$��Q�m����.�����`U�fJx� ��6���լZ�Z[��q4��"�����IԠw&��1�Yܹ���t4���� �ny��9K�]�nT��,��$�ܪb���!lg���I���K��I.��X}aΣ�]t�Uj5k�O�|j�8]��Y ���l֢F��B.!�Q\� �r� h��a�����[m��S5�&kVG6�A�F���޷��wppC��_
oZ��D~��[�r�r:/g(`}��d�R�YHX݃)�sHޠ�7��X�	Nd_��	Xi��*鮓��U|_@S]�p�i�X��lf_KK�	e�_}r�^'����.NizY����tA��L����P���J�ݠ��_|񏌺=��	�n�(�w��W��%�v��Q»�\�x�r�Ɯ�r/����D���F����$-/ui�(�����=W��S�7�P�"i�ؿ�iD�w4-Z�eዴ8���0Z���@<f���5�5���z���y���O�({IG��QF�Y��Z�:$zÎs��z��R�2i��N����4�e�O��|$8��dP�ϗ� �鰛���=.��UG����ͬ������7֭CK|Ǭ\�T��Ө�I|@�Ճн ��X0�Ci�z��}�Si�r�u		�i}DH�¬��tu>��Nb7��;J��>
4��U���(g���M�@U��뮦M;H�=�xT)��U�I���N�5��g~�͹����������� 
ѧ�fݐ�&���k��!��n$�Ԕ�=gS/v�a�!=x��k�'��C,.�a,B�?'u(/2~-K#{Cjϡ�%�P��a!8����dkmq"Y�T���E$H����fa��8#���K��0;�H�Q�_D�����
�W�6��u.Ӝ���`�ū�iC=,..U?B�]$��t%�'�ā����xG�m�=�~�����4�����+4Ɣ_pa��1�D uɏU�{���]�ru�W�h��N�d��><%�����d#��9.D���5�L����~��ɭR������@\n���.-QYtƓ���	H��\��K�DO��V"�sC��F�kC��׉U>B1�;�<V9�I�W����K�n�Z0�b�2]���7�@�*9����>d�� }Q��`nV*%J<��<�f�4K�HR�E��-��U�֙ۖ��(���n���1�Q�zW��\OV/$�얩C��Y�<�B���ɒ/P�U�{V�/�j��3���m3�@�b���Y=��a�=�؋�ub��ͩ����q�/���OH�"J@��,�� ��*�����v���)��	қ-�$xC����X����
F�xW�5�#F�N��J���=u��wmE��%E�����9��٦�9�V�Pî��N�#n��^��f^��0O@X�Q�Z(#(t�^�N��<�Z�v�M�b�dҊ�lp��pJ&�qT�o6�9^��j�ּ-����<
���>#��Ɖu�Wk�`-��3N˗�@ꛪ�=��=�_Ѱ���m�F� Z坼�N�[��L�������]�p�c��z�;4ZQC~���a��_t�K�MoU���Р/u��f���|��$q����5�|�i�� ~_l#��HZ� ��CJތ��uI�; M;ת7��Pi�KK�(���i�5^(��l*g��pA�l��
������Y0,�{E�g��H���xt�&סW����s�?��sP�Tآ\��i�i�q�Izx���)zĽ�ٞw>�4K�)�=y"#���ͷ�;��?a��ܻ-�>���5g^�]���c��2s�.�`]Q�����O���w#����4�"Y���In3Rm�B	��?��;���%k\���
��b��U1�\�yD$��-hh�@��X��1V�E6�NJ�Z4g����8PEGK�O�`��
�Z��x��ZG�R�/@�ײ�_s���A�$$��S�A�4tq���a::wh�5��(����ݐB�n���64w�إ]Z��T��l�c�Yj.In��N�}c�� .5ЏJW�Qe��r�-,��ٲ�6B&/�9����a�#�sם�������IY#���?���ډX��l�\�e`�r��S�����[i@�T��t���*�u�B^���"���8����6�&JSg� f2�=���d��C�.Z��:���v�ė��$/��'��>A��h��ڐ���+��DEʽ$ף&�@(0��RA��φ�Rc�U��)�YI[xI=�M>y����hٛA�H�D]���vGi*�`��t��D���H�j��
���6�Ϥ�1/\�xH���mY�� ��#+f�8���P'1<I`Jd��k� a�A8�QH)T�FT�)̲���������I%�1|R��j�r��JY}�>��&ە}K��-��0��j�K������FK�31_�:��(2;���Z_����}��h�(c�qnGG#{����}E_����{4F�^�a��m!ϻ�H���pqu���������k��]���S�x���=���=�C'�hP4{���3���R(s˾$px ��x��D���d:ќ ������P���a��g?��38d*,b����Y���N�75�q�
Nmޭ��Q���_X4����vE��cP��Y�cVn
H�2��(�A������IZ%�`�xoIj��W/	�Ҿ�MI+��̃����M!E��w��@�C�⺤��9?A%����������ҍf�'�`��~�j�X��v����8UJ�80T��B���w�8V5���H}�Gm�q%�
zz��_ɓ��^_$ƍ,����t�s�����F�kX�_6 �=B��|,5��w�A��}9�ء����N?�`��P���/�K�>�s�0뾋Wŧ�ɴU�?��`��;�!��m��U�Q2̌(叭>�0t��ǘ��Ag�[C"kѴ�����ER�%��S�V�!�m
ѵ������tt��I�h����0�e6�j)����	�O��Wz:d� ����-L����D/��3M; 7Ư�Ĥ���hX(ħՙ�v���M�!��h�-gUŞ� �"��~��50�|2�B�T�GOJ�T�Ubq�*��˴aKga�k,,S���0�Ah(�q�q4�H�?R#ҽ]��M�E��
6�b/0/TA�0�������˓�������U�Ϝ|o�C�`+A���|�/���/O�o���e>�k �El�3$�9sj�ys!�x�\A���B{���N�(���/*`[9��fx����J�4��^��F6 �p]�֓�b����D�L :���VC��a}�n�I��v�]���=����c+�͓��K)3ҁS�z�B1����-(�f��ӯ���P����K��x���n ;]swD_`�u�g���U��|��@b��,��D�Oj'��Y�=-�:8�ʡ�����R�c#����os��ݡu�!V�
Sr��a����Ԭ#mr�f�{^wa[�G�=��f�"�J����'�;��S�*��]��o�Z-+,��
�c�e�jV����
 �L#�2�����
�YOF	E*q�hh�0���ԓCpN1�J��w�?�o[��334���W�B:j�{�m���(�N�L�gUD��qB]�:
IA�D��)�&^�sv�� �,2P.�N��0��xs�t�S��9���m�����Sb����,`d�Z����=� 1�DYO�`|�9���@8��q�νܢAP�l�|�^jW�k�K�v��3�WKS��MF'���}��7c������u�2��v�����c�/��@N�h�v����ӂB�� �*#���'�f�;��qv�xϰ�D�ÐɏN�JZ���F����{{֪�E�W�&լ����x�u�C��H�GR�=qp*v��GV�N��k���!�#;5P_R"�gW�X�����i]v#䐧�5�7҈g�mW��%�8��b	-�b��fh�T4���)C:6�i"2[^�_2u�Q��X2 �v�6<��WKrʞ�~�cvT�4<�.c�Ի�V�o�l#��u�Y�?�G�咢T���k!���̆p;ٝ��y�b9�m�V�AX&Ͽ6�R1�5&��j*���<���S��G��%Q����$�N7xu���a�	���7�0�{Ns���B8J�g{C�:�]�>��b:?\$�H�s�&׵�^�٠���_箂a`<�x���8S�,�V�x7��l_���1����d!��w�%✰YY����0��1�����z�^��.ag<Zl ��q�z����$���1]쿸[N�(�㷵p� ���!ےB�-է6ʴ��j)]��.�<��[�T�;q{��׿G���x�E���.w���i�{��̅���L��I\|
�S����$�[�윢	�g7���l���O�m"%���HB�)>S9p_f=�R�j ;l�1�	�׏!�aX�X�D@5u4��POKb,e�r  �g�'S�^/��y膯��5�sԤZ�ܾܣb���"z^�׾,���u����F��0bIF��p�.8�1���ő�ʘ�u�{O������h���g=�ʹc���rX����Pu��eM~sZ�+��5���wa?�6�^��K��{�4�XmR�z0�A$�5�w�jf��|�8��KU�[�4ҽ��H����v�R&�T�ɣ�t>�'�B뀗�'֬�
����G�i���Y�5ʧ��V��Z�KJ3���)ka7�#�H?��0��+�,^Ks�[@�ؤ;�{ˁ�M[�n�	x!Q��˃B��hRk��bޞ��8�&��h�VF�le�w�k�Xk�ƾ��q��6U ��8�6�k�Y�.i�@^�qe�7��q��{��ٙ
�����m����%D�O�*�?�Y����1��#�f�hj6WYT�]�j����-<��k��Ri�x����6e$"̕�!e\��7tF��ԧ� Y^w�H����Zq�`Ev���P�A�r7j�Ͳ \��?���"��[̯�f)v��ߚ�x�Tݗ ����/Tf�h���VW2'�[x�d�iw�1��Z($��9*<�˿0����$d��)lӷ�/̳S�!�	�*O������\퇿�lW�q��w�3溌pcB��0�,2H�Xdkz���;�vٜ�to+49֯�C�c���.�r+�ӎ0ܦ��-��0����L�g��(G�?;8�kWVKY��R.��;g�E�����,�/1�tYI2�; ��}t�zu�z[IS�jg����Ӏ\���"8_Gw���!�2�VQ@jKo��] ���>(�������1 ̀r2ǳ���e�~ p��T���}BU��5K��� h�~�!l���i�|�w�&��<���R*l{�Y��d=.����T��P{K�K<v �Z��1r���.Yf�����ĵ���移_ZޗG�2��r����;p�7�$��?#��u퀗��p�?�=�@Oϡw!�l�x����+��@�&2�5PFc]ޤ/G?3�ԟ�q��r���:�����ƾS7g�~6.�Z���S���E���$��j�N�t��g��>�f�o6��&V@m�B/n7��� H�������<��zFU�Y��ľ0r�o���4���x[/`H�&��
}�~�����H��qu�����n*��sƋ�<��'��^�鶌�^4\�i��A���I�
|�����>U}��^���@Eb�=.%����B˛�_��q�	 =O�K�DG��of@�t7����z�̃���EY,�D��F$6�$��*d�����-W:HF4j5���$H�&v��FT�&������s�Ҁ�]ԙ�:��#�2�<<~W1�Y9'������j�5e��t�s���$~6J���2J���