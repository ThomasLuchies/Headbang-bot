��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q-��A��0��$LOJ���(�\�&�?S(���Y/���9;�g�875R�?����[����C�bl�]OT���V>b�`(�ZUO���_^'�>�F�
-�y������������ypڡ:l�����T+)G���r2 =��5BFn��'�1&�&��M�0��`�l�E��9ҭi�+���mbE$l6
ם��!���'�L��4w}^�E�f��}Ƙ�~���2��z��=�q�Oq��]���^�ZMY���
޸��Hn��	�E��L
M\�����yo��t�рf��^oG�BG�,l��	\Vn?�y�p��lr�Q$�(�<?z߬$p*Ɍb���L���m>&�\|̥��M�q��Q�UKwi�l����,A�n���ILL!`�i����t;��m9�ɉ)�pe��~C7��)�!�\X.~[�!�\.�Isq��S/��"�.T`j�=�bw���%^K,14���R5ݖ~J�Ĳ�=��B��J:�Z�Ol}S�(�tq2	,��i^���x�t ��v����}�&	Ac^"�;	$7"�j!jr�n�=,��e�]�C_��m�Dv��/���Vs���
S>�P��_����NZ�����>�a/�,}͈ ʸ���J� �����EH����y�lb�<S5҄O�Q��3[m]���s�1�5�6H��4��c�W.��]*���Q'寗���S4�ߗ�:�#��;�v|�_���u�kxV@i�c����"�9�ao�W���>�S��cA�p��\�C�R���Y(;0�����2��6J��ݾS��ኞ&��m�8d`̓{�^8\� �� ԰!� ��Su�e��hx�լ�Z�(bN����>^"(�)۾��>�Me��Ǣ*���=�$�%x�Ծ/�G����.s�@&��2��̊���9�1�&��T,�9.��Խ ������N]�E��A��h��,����?J���Ow���Rb��[��3֡����c�^SWR[���N���6�=���Ƚ2=g��A-����Rq��N�&@�Ҵ��|*��Z��K�=K���g82�~PZh��~�+sK���3��5S���>����c���>�6��3E����������~��cU=�� /�x��Q<f�x���"�c����?�'�a ���
5�`�>��;�`�`�fb(^f!��R�=OAD
]J(�D��_�Ͳ�sj��B��-�������S��i���l�^����D�ǃ���DL��8����-��r�W�SA��s!��,Z��&MO�q�"i�������R�f��%�|�X�Y�� �P�|�7/��1�=���iXn>�g���L���p&+����<N���XU������Z�xv����g%�#�4j����fߑgn��[-�ѭ��%g_/�$%�Υ�XSh���>�]�����q�[a�E��Ɛ����ܲ�ǹ�/3mV��V�N�)T��Y�DZ��q6>Sڷ��I�s��UI��p���M\� W	֛�~��k���_��m?��bF�cy���Fl�����/������ly2���d����Y�FW�
�A7��I\a���]�9�E������{�5�M�]��D���2����كw!����p�	ʡ��O���(���d$���:�^9P�ui6�
2�uTFj@1��UN�z[�7[�ur�}3�G,̯�'�?��Q��Չvu��U���0��{�e9>4��L�0�v<���W&��s�j��gP���Ǌ���!�2Ǩ�0C�M�a�q��������&�0�t���n?�T�B��?�'��E���4�34zY��I�J�oa}�gX�~ּ`��=�o�����hH�͞��t���n����S�)i�
��ore���lF0��v����4$[�� �+XS�z�1��eM��(f�fh�?��vy�KAo���*Zαa�	E�D�*P�_�E"��D9��j*(��4�f���[�Zq�LX�Eh�Ń��[�c����Ԧ��c\#����l��t�QW�H���1���YVݨ�f��$�~a��	~��Xh����Dv�ZR�����_I7fa Mc�e�	�8�W&L���cUA��1W�-h���K��m��T�����h�s��4M�ҙ���b�Jn�tn��8��Bh�:/��<\�$�cY��/���=�>���b*{�U��~La���u��;+$��\V0f?e�@�54&I�*0���-�����L#XM��{�CC�2l�L��hXR�"F���������_�K��IP�F��5Y����@a.����|
�IZ��m���OQ�RY0`쌲��1z֏�] 1����"i��m�3����"f��q�����h܊�2o6�l�����+*�0���y�0&�І5�>�bY��Ȕ�Ek4x`+�}�˧oU��m���ȟ�T��v@�S�۝�Z��*b麄�TDt�-.4`~S���P=̱<�3 ���pD�������٠F���n8r���YϹ�tl�����NRiu���/�%�i�#	.���ܷi2�h���	-5[lQ���A$k��JJ6$!���OwbW� *�Q� �Jm�|ඤ���$��d��9�7�9�Az݂%\ S*����Oc� ���)٤x��CWe[m������<>%]�Vgz�vxM$��o@��k�2(��a��!ɡ,�}Z���n�V�X0�uҊ���qsv��J;�174Ԕ����J�c\.4���J���V��r��+��~ZhIu��L�1Kr���lG��^��@RЇ-P��O��m&�c��Ϗ��6�k#m�_��	�ޯC�[՞e�L��!�.��vǺ���T�o�^2Yl�{xSN���)!�:~.v:b�%�B������7��L����>�S��p���w����/a=0�/�(��&r�܈�`�􅬖���;`\�8Fc��)d�'�HRN6�����d���/�����2`�]�Ӈ�r�`�C�~�L�.���)��;�T)ז�!yJH�`t��l^]V�G�.Tw�jf�\V��E �-�#�;�4)�-�4�v�h��9�%�28���++T40SѺm�}w�q Eq� t�=wH���;^�2�`fq!��Zʠ�,yR�,���y�lR�q/���t���)H��
@�gL��]�θr�̑��p�o���pG�4e�F L^i��-�>l#���.�U��S��Xk�:��^(g�)�XZ$l)Is�ש��t��W�8<_H+`����R����]?V顔;Ww ɹ��x CF���r�&Έ�"n���!�)��'|#�!7��!f~����͟�d�+w>��9��DÏ&�pP�R��u5�xQ�}x�?Y�-]x�>�/�_�4a�0(vH�|,��f�Z��G$�HL��K��?�'ۑ(�} M�I��{�r(�F�����@[j��%r�YbB/�g��z�f����F	��l����*���+'~�뼆���$}�-��f�"��%�7lDaPA�i�ja�!��׶,����5@Aܭ���\Yۢ��a���ſ`;�4�v�Zf��U��Z+~G�[�l�V������aʡ
Y]���+�Q"P��!�����RW��g�{�*�+L�*)N����a�V��v|������7���Z���9��q��*$ę5�Qέ���U�P��.�*�=���՝�v_�+�%��4:���0��p��s�ʹa�������u�wdg�zj��#��_��7��$Ew�����/(:���d\.��KV+�-џ��P?�\Z��#��B��c��0%r�y��|S��y��2��X�n���3������l�«r�i�6�,#�][׷�[�����L�C<��Ȑ�NI�u�C�!��~�S�l-59��AP���33�>+��uQ�Pęu`F�g�b�@rݪ������3�P��iL��[�J�cA�%�V��j��fR���_w<yɢ����ъ`n���Ͳp��*��*a�0�h�U���1�����
-}.51 Dg-]׿�Ӽo�h�x_boA��A��[�/S>h&���d�41�R�?۫��|^�5|����r�n�k��K�����=�OY6d.S��k�)1Gsӧ�_N̞�M�G�Re������;ǨF�`.��yE<d4�����T�$H���1��󂓐T�t�z�>w�B���c`3��&I�Nڸ#U�=��=���� �X�&�^����@�b���������6dN+�]��y[�KK8��@!��e[��d%���=o1W09`���k�b�'l�lc"�c�k�.d��w�'��v=�p6:�V5rn<�S�j!�:k�3R����^������P[V C;�fn�,k�8�1��d"8��H�������@U�o�{�����31P�-��������J?IĪ
$��|�y�������&�����«�����Β��R檿��s4\�G�.Bgj�=$h�pj��a�|^2vGS]�Sp��ϷI=eW|ͣ�цh�"�tN��Xκ.^�Y���	RxG���	���ˌ��J'(C-Y4�
��C�Ƕ[X�X�mf��x&�/ܢ�Ӵ���0���K�����\1x4��Fm�y��A����ZK�,�|F�ʢϊ���G���V���XmXWD�\R*2WY+����%�V��ܕF3��/��"d���f̽���-��[�~��^��4�8vCK�D�T�
T�h��Nl���9VTu��E����:���P�I�́q�`<���ڄV�w2�![���O�
�
3!	�k��a�L����r��ڊX������R�]ϯ�Dv�۱Dv����-���:ћ�*qѾHD�.�'�:G��R\T��&?׷����x?XC&6j�qf����e�<?�����g��~A����g���o�=���;����Ϯ���p������~u�*��<,�.��z�J�q����<�n�,�zUm�6���c%�1���=,3�/�1�b�T��j�.#�'[�� �tx�cZ���Gk��D�}��Qf+��!߈`���Ĉ1쭨w+�v+;��{�f� �Y��Eh{�
�j;B�+�\� ��q����/�3g��ud͍��Q�6�,ً�p��#���7-�S�� ?�V��"�-��Y]r�7y��֣�x$��Jr/#'E��P��p�H�a]�pO�K�_YV[*���]NԻx/9�ZI�H��:r{w��"��-V�5�z`�H�r���I���ch���;{�1э،҃hb
� _�0����V��P{f���RUo[������j^��L��V'S�fU�䎟�M�8�����	P��Q���Pq�ؘ�v�j��x� {�7L���Rs���Fh���z�2R��$c��y��[��o��5��8�� ��Ü�3�X�v�ȩQcg�� ܃���ҔTG�Q��M��J'&`���x	�Y�g��|qF��)<��G���rL�80p��,��<qr;9�7���73�� }H$Db��
�Խ=T�FϷ�(�kA~�ϒ}0S:���W C�g��ֺ��� R��N+�{9�̡m��)�Kp�j�/�f��^vMޖt`z���xQ[t�!��lI�4'��m\�0E`��e���){x��é��PMe����:�p�xc�2�1�\嫒��=ٶ6(<�ϛZ/���k>�����<P��ǥ�ꐄ�6���K����ڮa��<�h��?|�\$ٷ�Y"�2�J\8Mr��p�d�3��b��Ӈۈ�JQ�Q
���qR� !&�C�=ob��*�,��c�!)x�B�wJ�)C�Usn5F�(�w��Q��[8P���s�n\�꠆(Y�;wp.4�m��;`+G�k��-�?���2(���L�L�0�����ƭ�ǿ���x�����L��I�_���U��<魘�<�G׋��[��i���[���,�-��B�S����v����-3�U�dr�~��)�/���vc��v]� �lJ�`�,�c�EB�ͰŬ���l[�p�&f�i�����2�C��B�Wcf�N<���LH�Y����ROwU��p��q���m�x/�RyR�ʰ�@ެ�i�n��F��jkw엙uAs�T&�;û[�e�����^��~S2"��~�~����^��m���n�O���H���r���@�P2�	I�r�f��(���Ī3o$�],���k�[�����$�g4e���j�*A~��VL���jM����Ԕxx��!�|�(h���g��uj��؈m2�����`��7����H� Px�-GU���Np]�(>�I�s辴V����o㖰hH#�`&%H�y�@-������6�VȊ��G� HC��Ky���[G��F_��g�>��Ȑ/�@�����70 ������(F�ȣ3�w�i�!���.�D��h-@������F&��O��fm����R����quH��8�����ϊvt[D��]-��z����+��-D^ƙL��sRS�+3j�"%V�Ct2@yI�LH|U>͂�n�y��="��VӞd��GA�[���؈�٘J>��Gt������m\�\\�D4,3���r���[A�U��*�q��\���Q�%Y�(+�h���)�l���~��-mT#s3B)3��Pv���q��l$���c$��F�7۲@F���0�@eҺ�0Ӛ�[�_�<��~[�|�C�D=|��ߣtF͞,�W%3�VԞF�j�z8$��&�x��9V�k�ɰӕ�(u�0N\
wO�k�LW~��yVf��m��o�TS�T�[�O��Όq�LC+*5��3�+������0�
R�D�k��%��b�HF͵������t���{m8��,.m V ����+�߂�z�'?�I��R�|J@L�uЊv�0�4���+�*�����U�!�;�}M�r���G	��JA��g�xeu'����̫�ه����πlQ1�e	�3E�P�U�T����(��~��|����9���e4���k&�_�³U���[�Sr'ꌶ]D���,tǵ����} ;,g�Sd2� zp�h��j�	�=���g�)�@�3�fI��q�- ��EF�!��� ���'q���2���x*A�](��UA�#�@�WϾ}����!V���Ǐ���b�M��_/F���-�%��UW_Er�4�#\���X�v/e��,����O�P��A������Ʃ#� ����O��G��f_�%���k�'�,�N� ;3.(:�}86�����fdb^��Dn-4��87[2��4������ʹ����?xã��y���c���[+�L�o�y���)����֌�sz�D/��K,�Բ�n_9O�����g\�]�U��f>
D}y�Y���n�p��p+g�_�0�ȍ�5)��|�Pݴ]L�*I&�u�Ogw�0��T< |S:?�]�,๱S$��IsA{xSG7"�S�c�|^���t���!D��K�-�|.׍� ���8Nh�2���䠸P?@*��XSE�^c|�z�5HV(nJ�?�����Ora����T���<Y�=��l2\F�Q3^,���p�f_�p�����SZ^�)@���Mvl�ƽ���2����%�μ��tf4li�)��ʄ�#$D�>�&�$�X���# ���d���+(�}<����8Y���|�9p[[��)~�?�y�Gb��{�f���Q�=���l��䘵×?~�D���sw\����r�7e�9{S7b0���T|]U�į��g2��nu��c�f������3$+�)@��>����2\�3w�}~|�S��q�D��������tgE��
���W��&4`�lA�|G:ȗ���{�����u��sYr�^S:w��A��hf���	���/�"EV�Y�FW�k�7��%<���l�3�V
�n�m#�˵U�lt��+�ut�V�z�ͥjb���X�!M˪L�4�D勈0k���/� �x��ZC��l�+2/Ԙ����b�_#��Ԣ=�$��}m��x�H�v��v{_����E��hs������5B�<+[+�ȫ7���6�x��9O��Jdŉ��JZ�pw1��V��&�Jퟲ腡���^׾]?�s�5Ϝ�����HLP(u}�$~���#M��B�6K�R�goYū&�,1UH"c�hG�yW�VA�*����n`R��}L�P�\��p'����e���_���b��V�
�mH�3�^�(3?����"�"��{�R�9W�$����
����f�%+>8���X_�6�lt�͟���M���Z��`�a詅������- NO�r����ڣ�Zo�E�+7A�jt�m�<O�#�I�~mk���!���oJ)���7՞Hɋ�С���O�ۄ;z���M����Le��~�`u�H�c�����_R<#��B���3#��vC�{騖�q{�*���ߋ*7��������!;qi��؍�qn�$���KZ7Y�ST��9>T�W���au��P�?�A̓2�'c�!Jz�P\0-�ȳQ&�j)�u�F�ӊ:n}b��k�7���.}'��P�'|��z��L=��M��qe�NS��F�cm�%���{����{���g��0j�D]��e��@�9��+���.�]�|�����p��B�[JK��(Z��mN�K,��$`�
y8~��^/8B�u-(��M3�H�@�o�6�	�
�H��ܶӧTD�$l~M-%��/?���l"'�ж�F���{ DO�h'�.����V���	�����Z��G���C�l`.=��H����gʾ@�&�� H��Fq�2�b���5l�]� ���M�{0���"rl)H#��C�O(��d-���K�e�����]��<�a��!�,r����*��7 ښe��|'o��Q�H�趯�#�3�\�^��7�i��<���_i���z���I��v���8C�
Һ�.��.�ի'�������3WFV��TҮ��ng�M�	�cw����r���� +�f
I�s�Q�ڬ�,f���q[�Ϊ_K�|�N���k���X:�b�m"ݛ���p���9�B����R{S������ߤ�3���/m��v�a/�!V4|�#�M9�`�	p�Fp�������B5��&���wd$=8��g��������� Xȩr�Q��E��	����V�����+�N��b�{ˮ�a������i�q�e]���9�f��Wɢ������<��s�����y�r����PX��Q�@d�z�J��;�rk1x+yY�;REM2�&��zĨ�O���ߊ���R���R�[�L��"nH���g|��g�*��xE�[>�R�d)R�����U�퀩��_<�5�����ON�!g�=�t��ސ�t�d-Ù�#Ҿۚ�3#����r&�n����C�wx��A$�c0 fy�ѷx�k��	t�B�K��>4�?����Yy�g��)[8삙�;��1n�vw'�_���_5dE�4�ϝ]>&��3�,UC5��i���w��}�!��T5Rm/�/�G�'�\����؈C��?�/}I��i�49�b����u�G����!i�÷5?O��h-�X?�����k@��l��MD��o�%v܉��c��=�N4�W	����-V�:;A��y�J)+�=���]��Q�6��&�=�g��H`4���n×o0�#8�,�rܼ_�ss�lS��_*^L�"�Ru ��=����0dj�Y텞~Q�:����X�J�{E��?��QV�:(�!<Hz�x�럪p6di��i��r�:���H�����3��9��f���7�ԁ�T6L��/o��R��ڐ�'(��"���*��'k�;°�,k�8H^w��mRd��1|����s����|ڝ< 8,��&�.�� �E��4�*�}�6��L��@�SʶPD++� ��V���g!�����+GKo����-mW�6�x�뜅2�����q�$5n�$�C��$<!O��}V����L^�%{͠=9���4K���w���� ��	~��������_
��Ñ�a"Y�� �P���ׇ��� "�rS�}�=�G�y[Ô�۰���O �t��i8ۓ�
|����w�gc8.l���(lD!$IWl/��=��v�lG�]}�������p�*�-c��;���"�N��1��� ��FPG��42�HH�&�V�D{��4��Uh��v;�yiZ=_aX8��3�,&`��e	�;��ƊHr����q&�i�̞�$��}�ID���@<�y(b�f����$�	�@(��Ԝ0���g���%�~ ��c�����ҹg��qL�D��3�d|Cx�{٥��љT`H02? ���{�.bp8.�w�kL����ʶ8��6ϩ��y� �/�V� :��8Ԯ(\�!��[)��,�����qS^����b@�K� ��i�A�k���r:�ڟ89m��e8o�8�d� f�v�f��HI��#��WC���=���<@��Z�ȟ�;5�
� ���+���n�_dJSJu�6�T�V�#��0���9�A���Wf{a^��k�Q��t��X�����Fy{�����="� gD8ݕ��M��6�]�p�{"UQ���ũ�߳��;���??(�pV�f���x����?�+��z�pE#�q����@�l�٫Z;�n9��'�/�kג�8aMb�~��{�M��_xRS^�_����[����h����wb��8��&�8��)����$Ruq�-�"G�(w4�Tg
qM�Ya�����tB�9~n/�s#������-�����n�F�y���Z�3�@��a����S��4�PsC��3p�B�9�dp̔�S�]���Pyya}7KѶp���٣�gl�u��g5�/'�莣�î���ߑ����aX�U�/(��8����c�L�!�.Z���=�^�z���4"���I���3�7�����m�m�Ȥ3�_��{(솥N�к����T�j�Y��7Lj�0n�%q�$����%�sFV�^�Uj�@<���uw٠��=��ˮ�F�vYV�@���Fڧl���h��8e¢��sKh�e[��ȗ9gs ��J�9��o�N�#��V~�^*��f���AR�PKL��g�d�(������ZmB7��{����wE@+L�y�&�U(��,�Җ��;��3(A�*�����kȜ7��O/!�i�������0��z�D��8�rc<z��"� ːB{�O۳��4�����2l䙶ݑ����T�������n��t��Ҕ}��7�#�.|�J����*��X�%B�%���6�(fdG8՜ܳ(��`z �<�pا�@}�Fep��kʄl?G�~�gh�@W�B������A=k���[����a���)�2J�[���q�t>�X�������X����͹G0T��e8F���7�3�]�V:M�ς\�����槠�Kg�{�3p!S�'k�����ϋ?ƕ��
����
$W%���4���`~K�GPiSTUe����'BcA�B)��xK��J�i����X�Z�R���|y]�A���}�˜5U��l<����K[�q	"����N�A� %(Ҙ��^7�1�Q��@�Zz���3�L7�0N,�*ѣ]j=.b��+~�O�_4Fe6�
�t[;`8�ѣA���і������d��)��G�����ʤխ�e�Ճ�l�?@��O	�}�r������ճq�Gr'��ᑱ`�$}W��̍�P�J��3��n;���@�@r�w^5,2-gF.譚]2�O(��H�*zC7�W��Y�Y9���oԭ~*�EF#��ܓǦ����\%?h6d���E��!�/�65��<�Z��<`�#m_.�eɒJ�XKO��y�����I���QA��N�L@ߌk�)ڸ�nX�h>T_V���襍y�`:<�7p�N������>��C;��z�����G�~�_,�4�aW�N�������gR�SӞ$iP������M(i	�$SPFؤ}!'�TU����(�/����"�N�5���#:��*��DN�QM��X
�4����������s��EC�s��$^���r�~"R�A�>�i-a�3��8��|C���/�����v�7ˆC}:)	�6��1�StN3���u��nWByK{��-�Z�m����V%9e�uѯ���q���Ďfo�%�X��\Uq3�>�$�#ߗ6�=�0�6�^�!gf"�[L�~]):諆LjP]�2�"���W�{p��c���\r��fa�o�����b{�f���p�f�q.�j���O����`}Cd���4�.��F�[��g!lٱ1ߋ��A[+q!�d ���9q'���iPE���"�a���z���0�v�kfd!���|��ܾM &�Ix�D���� ��8��+����=DJ&m�6�L��л6��p�N��;t���GJ�d	�%�hZu`y]C/U��8�]���5��g1�P5���VR��|vI���7+��9�3G폧�$������$�E�L�ǡ\�0NAiC���o��}���*`����Nc�yT=U)�6�'=�H<�S��UX���\����%D�C�-��~�/��d�s�ɜ�H�T�؆�yI/w�$ꑵx�d<�0Z]* �����_��l=��3��4�bg{��T��~®�@[�7��iD�Y���V�%�e�䊀�	FQ��r�OWʥs�NL:f�#Z��0��A۩�wF�m��0f����q�Bs6�i�o��Y|/�@�>��]J�l\����<�� B^[��,�E̅h�M=[�wt���b�XY7�wzZ�/ꨫqE.�"�_d�� ��!˭�"T^��c�Z��:�	y�DC�0i�9��{��:-0ެ�O媪ElN����,�������Ey�#�-�չ�g�����ϙ;><mx����/A0���Fd��׹�8w�/e {K�BPY6CCx��ޮ��.ٟ�v���B~k���d�N}q�Wz�,Bƽ�呸8LƠ�9�A��;��0Ί�k�ٚ���5,��AY�*��SI��X����kYsP�׷P)$��T�ᤂ������9Jm$�����s�.�]$&������S�h����K(B1�ɮ���6�;�߫k�]�;�=�r��;��%�����rUl@�e0�n�lX*�\\�N��A
��j�1tX��x�Ԋ	�(��8�n{Ӝ�� �,V�ܸ�q�:�ӫ ��<�2���G�y�Ɖ�Z��:ЯC��A�(K�y#w��`KG�g;xq�Z=�#tP�$X�ˬg7!���WlA��k*�B��q�Z(չ����*d!�]jXѿ\p� 0#RD�i��'��|7�:|Ĳ��K�]�/��&�=�y����B���W�$੖�K>|3Ex4�-�
�WPQ��>Ο,�I�>�r���*�ʝ�x��N�Z�6���$C��"hn'�\X�~!����U�c�>��_��-����)?9M֓Rꒊ��^����}��.�c����MR�/1K�&!�����h�´^6z�:dΒ/�7��+��e���x6�*�9z�ZF�zZ�x��^x�@��#�#��,(���|�����;l���o+Kɽa���2?����z�X}ʌ;�Y����7W�%٠}���GYj5N�^Z�m���J����}�)����1�&�����?�/�B��|�Ir�>F1�y.l���k9��F���W#����(5����@�4�\1���	�`� =3��3J����C�@Z������gTpj����E�Uh�0D})}�M�z�B$�I�#у�0��� �� ` 3Im��r͈|��@BQSLh+�tR�Ґ�v0oބ�y�Թ��/T�)��zt����'�r�M���$��hE���FJ˩�Eb�)1:��% �/��7�^���c��1�:y�
�fB=y�d"���}����iY��٢e[��&�������q�Y���¾��I����얝T«PhG�a\�E���F�F��47���DLJ�,�F�Ԑ����`����d��$1S޶�#�;~�E F������MS/�b6��8�)�,O�ǟ��� �i$���LVj�o�DRR�&�1#�!.^��
h�m�<�i:v��wL���`�P#����6H�e�"���g'��2)_j�$�'���K��9|��@�7j��$t�8z]�Eu�(�o+V���9ɦ�k��6B���߸b��EmK���)F@�e9�p�+�y1�5���؝�6��[�p�J?>/ȏY%����D~�.	Z�/��|h����*���.9���1�gJi����K�,���oY���C�'�����Y	�?B��Ɛ6��JT�ǖ�UL#�'����┧�b�S��H�M��&���i<<��7�:����p��7�{*СP��I�F��Mh	BPJ�D��.��YT��`�w�?h�h�K���3򫦸5�cg'�l�0Bⳮ�nsZj�����?Z�C�&��p���\�0��S��=�ԉw�Dd	��֤�� ��1�g>'���O�O�\�^B䙀�A�q�rRY���%��!,��@��}�ie��#S�N���Ub\�k�b�ZJ�������=0j-��H���� ��¾��{����_X��%�9afG��8��iu�	�M*���=z���oa���E�6M}�� W	@&�E�I�PCd.���)�'٭Ĥ��]~���gV�A�;)����p5��*h���=.�˦��-O���,�s�D:¼� ���
v��M��)ޫ�-�t(U�*���0n��,�����=eW�� f���98O�VZ�86�}�BoH�;SF��]����E;%�$��}� �kˎ�����p����2v���������7*+pH2����;E�Ԙy�R�ݳ�є���o�p>�:�Α���O&���@e�}�d��}a@%*�iP���x���}܅��?Èq*={pvp �j��Q��$/��[p#�v<�E��q�o��H>�Ob#m(t��Jv�J\tTpT��M�?��x�pS"<��R�U����!艏H�`�Ko���5��b�D��u�ʅT:L���&4��[�e���$�~�?𽸦^$D`K���y��^�O��M�Gl���^� z�ԡYZPM��3Ŧ��7E���K���0����,;¬|&n��2�#�L7]a�I�p���<:��4[�W�L��Jυ;߿�Mw�?�:$l��ł�W��*�擸��agYx��> �nΚ�o"נ���PY��ʟ|��sB^
�֭��󯧴����͔�! �+ة��#�(X��������GjpF h"JWל@rb��:8��/�"F97}��T2�+ (�����b�4={e6e��.AE����9�����M�����R�l���e�7��@$#�u��&�A?���*A�s��1Yg�����i��Ե���1�Õ�JMs�-I�m����?�1��S@Z�=�G��%$l�������r����d��UaH��=�>���1���UAѨ��TN��8M|�k`ojP�瑡ؖ�"�������\�@AHK�쮔Yn��[ئ~|_˽0���5�x��ٺ�Xc.�T�z���97�E�a�p�)U)��&�$�c4�=�kun�BMo4qQ�����39d��)Pz@�?��]RY��u0Vß�,.H47p^߆CW�	U���ΆO��\�J��L�*��n�Ge$P��D��u�+�+�p�J��|��-X`�1=�K��I�T��X�.���;'���vpD� ���n`���_H�j��p��kkRU��*�9.(bB(#�\D��_^�O�r�_M9��g�R��Q�����iª�&�-�V�y�І��dq,���b��̴S�^�u���]��-,�=^��W��;�x�A���D���G�E����n�H��Z��x���P�Q���8�'��^M#PW%Vgf�����|��R�y�Ö°M,-�p�k>��a9��)#�?3����}>=I�}3&A��"c���2KV������jS(R�i@����{��`M<i8���Hc�1}�&7��n5�˄��p`�}S�+�xc��L�o
�G��u	?H�Ƈ��MȐ3<|�r�;C��U:N'���0�gI����������yg����j�3����W�����B� 6��o҄b
PE�P 9���Ljo�c��S�"ix�t���) �e�')���|�{�G��[V�Կ#��!٠�P����~Rε��SY���&1�9hϮ�"�I|@�:�I��p����Z�H���1O&�厳��CB��4Ļ���a�6"n*��@��Xo���ڳ�+��t��E��+�D�/BX<v2��O'�KV����J~R��Juz�8;�bFbV&B�G��K��Y��4)e�/�c)Se�Ӧ���R,��&A���A.=K�F��e~=��Ή�ÀO��E�9�[�Cm�����|��DQ:�Wߘ�Ql��}|ߣy?� �=�����FWVc�m�w �8��f�4)Gk�Dq�P��Ǔ|0�`�+�J�%�G��$��T>!V[��� S8�7֟�/�9�<�+I��[	i���H����;�0Cq9�^{�d695�����n���`"�U��� E���g��W��R_�Z.ш��i�H:!s1���M��,W������/L�W���9Ed8W��F8�懯Cϴ�Ů�}/[���Ø��W
lh��K	0�"��������<�w��`�f~Р�듹�ھ��%��7䎐{�\�Vo��+�.Ef�}b��R�h���[n8�oo��v��v͖m֋t�ת�pڴ7��y;��h�l<^�x�ҙ�#�1�6�l�������k�Bjd��J]t1wEڴ�~���ĩ2��x/��ޑ0�T'�1�R��n�U����������+k��\�e���`+��'F���A����U��:��U!t�h��U�L)�����)�v�+��E�2W#z��(�9�rr	m�C���䎧����j�V��i���� �i΄H��8=9�t�-��o���8R������o����Q8�]�������5UZZ�>Ԓō�y�l�m�и=��_ˈK���y�f"|uh;�������(��ۤ��[��b�l7�|�i <nf�b��	{�:0�c�����ej�yү�e�*�!-|�܆
�H�%�X���U����jR%M�
����D�E��9�h�&&�%)��"�#��'�D�M�)Xn(���uM}�x8�MN���2���������w�E�!e+.iS��@������<�g���w���`��0���%O���%ӭ���AŁ3����n�m<���̂)Ў���9�w�=%��5a�qII�WB�̈Oۯ��!�.,�ˣ]��Y7S�\݋�+�^2�ǑI@<(9W�C2�}�ZQ��� �n$�X�g���3u��L�
��\�o[��D�O�u��״:8�N�9&4%�#�	��s�*��|$�A�ּ��8I�6�"�HwkK�1.{��U5t	3���&�������t�.�T4��Uv�{>���!���LAGc�lf�A�<M�:���!���{`�W$�*z�1�6D%���vVJ��_��((���}������	}�9	�؜w�h�ǔ�`�t���޻���w�	�"���ag�/�K/ƞPy�̫�e�V�Ej�FC��m+��5d��Ve>�W�^6�$��ò�p@�W!�m�]��ި��*^rU�-P^�	�n��!��?�W�mVbJ��Uk��Ȋ~��UCqi"��+�2@�;�$4��m�0m�DD�q��ŁV5qNC]y�\@$k��ů<��g[��x�o��s,$�Y7	31|Q(�����EP����AF��#���wi8�y,��[2f1�|�^B-�i�s�8���A�R\���،ف�'�������u@�=�?d�)4DFw�c�Q�
v�lk'��i�ݳ��a���O90֦�t�`�r¶]m�.�!Xf����r�P��`���O:/�%�5�(v�¿����1,��m�芦��Az+��/ܦ��)$�;��������L��a����AS�iU9��V����E�s�J�f��~�k�}�8A��״�G�݋�f-
��X�"��Mp��]��e�q� we���-u@������a>�y��|4&�.�ڽ��U��!@cN���B�˄�������{�F�FO=�d<Xb�.�h�[��/bqC�A��pnqwڭ(s�=~���l�s(�"���0���$�������,��)d�� ���i  �׬eO��"���`��*��$��6X{+(BU!�����dON��
譛�փF;f,����8������ȗ`n}�1E0�b|��κ*�;��R�X�!��7x(�}�>AZ�\�\Ќ���$���lmB�#S�m�,�m�k�wf��I�3������C���.#���������� �?_QwN�X[I�պ5�!* �F�XjT�� 4�9�����d~�
��|��'[�>�TF�&�	�x���|�����ʺ�(^$d���H�~H=M�u�u�����Q�"Y���m}Wk���G�p�_"�#����I�P����w�MZ�a��@Aɝ��
"\c)�k/��oﳍ�Է73���� Kq�:|.���:gxQbry�-{�*��K�+�О>��91�K�AI�F��J��po�����S�x�M�q'�F)��S�ccx:�l�Da?�㣊紈|��n��m�hl���a\0�Ƅ(�a�M�3�|��xyS�U P���6D��S��4:�/=��E�Jך�)��;��5	VU�b���>��6�L��Q���"��'���W	a�3�!� 'z���66]�]��Ù����r�����H�����1F�lEK٥-1`D��D��w�	qVo���T8��'�LR�d�C��˵�a.���5F�_S��ըX�Z.4R
�ᜧ�:f�2�m��4F�Ӝ�����?$r9gE:[�����x�W��U�R���ALDts��9`
c��LX
�z��[zpj�L~�=�&:&r�
�����l�ݚ�1�#(����q��Wb���L}
�a)�+�������/U�ڃ����UmI�s�Y�~����G���j�_FF��}&�F/�_� ��:^���#�Ȍ�>=r�IVGߥ�3n�6�,vPȾڒ�ީ�g0;�:��[��ܒ�=/}�=��4q.B��(E�U(K�p�l2K<"zJR�l7̷�6��I۫��^� �QBʺĤX��w���]�p�.�3-u�U�f�-G�c����
�g\�W1�2�uH��>?�oM�Y��G$~HW�J��޹	˻�@M&v��)���l����UBZ�ɝ���v�5NIq�o�{����sb��P���p��,�J�/�70�d� ��2v��b.=�H�:OĬL���F)j����-�#d���O�������\0�[>��o�����θS4\�;MS!��]9�-Ӑ����1��m`0d;�p-7;(F��m����0�t�����o
+g��#�|��i���|��HR��H��G���`0�$��Q}tA�ٌ�.�}�Z�J.�U\t
��d�U*Su�m2��mȁn��e���Uwn�5���b����:������
ѣ��8r���p�IP$6��2rT���7B/9��`m_>��߁��PI���jTV�8�"j	��T�ENq��mը��j�O�3W��'�F�d��\��:���i��]�:�����Im���#�`B��x� CS~8N��f�ڊ���U	ُɡr�b(�;!�n��7@��0tN�]0�W3������((�7�/����Z_�@��~ =N�A�j�����2�i@���G�)��B	�t_�	��]<͞\Wr��
�M�Q�O�������9tU9E�ܖg+�1fLg�C�uS���5���bܭ3�[�K����YŊH���4p7�ü�#: 'w�c�1��@'��Dd�!
l����p��@��@G���q[3`_,�|�k���\��,�JČ�ĵ���`U�Ni9pK4d�U̾/ʔ�>��p;��S|��i�0< y��j���Q5�x��ܑF�m�ґ0�I�8X�ɀ�Wγ2�w��z��V��uh1 4���i�w�|�ܷ�r�r�]��]��\L�^&o��=�KL�$44+�F���e� ���A���7���s�b�푶�m��ް,?ie���'�ڌ��&��Nl�]��2_34��:_띝ON�}U|z�z4d*w��EOc�儽�ebr+s���2}`�5�F�������?(�/�ozQŝ�2��������ɘ*��`�桫
�Y`�Յ��JQ-�W�����3��)��|�����jgVF����F;���Jo�Ho�%*h'w�h� E�с��X��X��.�=���ֆU�N�?ְ�-�WJ��w�M��	������<T��`W �|��
XѢ���CF�02FN&�׫&�#&ɻI#�P��=���Ş�ǿ̽��<$�sވ[��rv����V:�g���� �EP���ȗ��NcrVL��������a�����s4_�׫5�J'�F,�$|_��;4s�}@O/�
��R�,ґ`����J���9"Xuې��֖�o���AS q�����k��s>b�TttPh�����t�Qz�B��L��r��8��18�"~��P�Bx7+|$�I���l�Ϋ��)=���TaPBla[8�0i��M]����>���6�w�s94���Ł������ 4�	�ܳ[VOpI!p8����𢃤[�������������$���c��c�2��ԇRR��:�(����'�i��x�`*@��΍���,�0�?Y6ܳ�!���|�Sg�`d��J�66)"3����a���r��9��Ӛ�����1J���H���s��9D	�9�|�{5X	?�z�rq�vq��D�A�v��w{��f��Wc�n. u�W%�k���#A�u�5w���k�Z�/������2-��yy��"K��{�ߢ���� ebD]d���t �b���X�	��S���K�/$���$�6R�^���&VO��q�!�	Fzq�+c%r%x������Zu�@��7_5���ځ��2�2P��� ۸(�$�-N�T�@�_Iن^�.�[N���TGѻy9�g@����E�>���۝�+�S��� X,�y��(��s_��:���~�X�S��rA��͚aIu�VPy!H�P���[����ђ�Ml^ƀ��HD[�}�]C.�â��-\�D�N�˕٤��^ &_`�:~N7�}9�Yg�ڿ.����G3(6D�]��S�l���_���u���U��v��⫸ҽo���Y'C�oR�H{��iP}�b�E��3���&d�x"�SsBYU@[juo��ģԐ�o��J\|�]0@��e�H�ټu����)�1o���f6I;M�@|���D�0���R!��'�'m����!�w�gh[r�O|�V�f�g.IHP����Z"�BFf(�������Z˻��E���PFfM�-�ဒ`|� �T��0�yH��4�X����m�������Za�����EB}Hi&�BOZ�)Sy�:�#,.�q��,zO{Q�����ڡj�.iњ½����*kC�N^K��a����r3��$w�I	k\�a�F�Ň��z�wQ.��4��< �E5g�.ރK@G��_��"�����UM}԰g�'�svJμmN��U�0C]���aI���0�(������̅H'G.2b<�������[�_���E�Ly�'"?ږz��rDJG��R˄�)6�*ZU���$b����_�$��$������L�])�C���'P�e�2m���� �<�ml��4��P ��������I��hKG�K#��q�.�et[��h��?� `DF��7-�.
=+�ݮS���m����b��O��l t�F]�@����x"Wr[5S���A!��� �
yU����� �z� ��b;:�;����L���y��$� �1�ċ�_�\�M���j0K���|�mѺ#�N��M;���.O%K��]rA=x�(�%�X�%�:d�u57 x��4�O��̓��'�z��=��Sw���Qެ�͋���[ьZJ��V#�|b<'�5��
�����><F�(	�#�p��R�~�j�*
�Pm��İ��H�C�^S+��e �q�Y�{���bd�x\nI�b9�j��_�|�#�H���z@O���t�����^����E-�n;*,FZI6;�8�2Q$a�J������'��;i5^���+~M^)y����;���cN�BI����˙þ���'?ݕ�����D<��P�A?+���C�ںھm��Id�9� [�~ti.8��Kv��>+t�9E{CX^'�K���B{lgb��32����i�Df�v�>�1��t;������؆~j�9:,9^e��-�K9�%�r��)i���2Z��� �ֆX?���p^�(����7 �S��Ʉ�rϏ�S��aD5��o��ƻ�����2�4�A�W�?�v[jqJ��u�Ֆ!���K"��z��+LU���O2��y�Tq��U9!�.ԇ\Z[:k�\����T�7���������;1�F��,­(�O|7�[�U��S��ݻG�O���Jx���0��<�9�'G�.�R︖��� !���5ps�v��c5��^��U�0��7AW%�(.bHڝ�cf���=Tk��BE�i�}=:w����Ŏӎ���fr�ٻm;j�ι_�l��"q�'!s��0cBX�"=��f}��z���*���'9�(���m�/2	�p�p����pr�:�r���w�|"�bLB�$�o*�:�R�]��A@7�4�ರ�pJ7��n�$���4��4��~V�m�y�:�_K|y/a����[;-{���[��#��3|�tq:�>a�i���&!ؚ�Z��cӶsH�V�x]�{����ƈ���0�����[ ����� �����wՈ�k��7�ϑܭyq2w.3<������ٻ�`p8Ur�\���iz* �A\����[#��/0a��%E��|���]!��ݧ�L�c
u�����z��"l��Da�ޯ���7��d�����6��_�/�02���\�҈i7Q�+<�ea��@Q�Ǜ~��ؚ�=v�g���L�)�G������M� �B~Uxu�c@�ט��:N���B�����l�H| �Pp�����ꢝ�������S�QTv�jF�N���E�3����%�p��T!�L�����@�&�e����(��
F����@?$V]�c�nm�D��&اa�PC�g�e[�&�QC��"0�D�(r�)gr[2�
�K���T^��^��9��_�1�"�}I�g��v�k�g�G�G�ޫ�*�?���B�Cw�C͘k�FK�(�.�^����+��^�F� =�<�����V�'��.�����fֽ?nԗ�,�l�|-��	����`W��Z��
M�N���GD��MD�"�YI��c3�)�A�Kc�R�-/g3S�ʾG/PM+Ou�J�����A�\�q9A�p�.��Ad��@*���c�ԛ^��AI���З.��=U�5W�Ͽ�lT���3@KdM�2�˔D�/BA��;0�n��;o����3�Yá�4��8�%K�^u.a\զf�1�F��R`�1��\d���� }&"x�?���垠kgr�~�G.=�?t�a#�`����햙�k�	��&kU(eL���ᦌ-�vԾ�?߱��H��y�	�ɖ�R���ҧ�Wx�}�1�t�!dp�T:�cჸZcU|�e�]=�dGQ�@)�X joE_������H��2vBLM�A^���T�߶y����x�_�G����l�~����)�r�)M]��W@Q��@�jZBD���5ˋ� ���Ѽ9����%L�M�k��j�� e�#y��y����UK�%?�ocJ?HٱÕW�}��E>qnZ�J�`������nߨ��e)ՁX��a��l�8���o���tH�X�1�r�w�l�	���f���������F=kOv���G9���h��SI�s�,s�	����'s�O,]�/Oƞ���gZ�x�6ރ��C�1��<Pu�ϵ?���XKq����u��Ğ�.�	�׮������?�,�e�aH'$d��w�(�;,w!� �!��'�"���n�;ƚS����Y���~]>�p(����,��ﱕT���9��t��>��&6C�<��((Fb��t_S�I"X��fDXey���)G��&�A�Y�Vo �uH	]��� �������K�޴�0��;���p8B'�:^CX)���f�<%���CN����s�����A#�#"��kj�| �6�&r���t�%����,4j��ڈ	�5Z�� ct��`ԂB�i)k}IP=�-@l���s?�COb�����nN�hsD����ҫ�Qkc�'�o���l0���Hٰ���_� L���F�=	�U&Q~ ����4�[���;
���ۛ�M3}�/&��+4��$)xb���Q\x�v����$.��a���K
?R��Uc���́'�h�n:NA��@dپ�o��+.�zP�׬�_{��&��\jb(](�8n���sA�c�$7�X��i�����B���䐭5#U�C��΄���	o=��K菓n!л�2���:�0'	�mAj�σ�J"�%�P>S��9U�Q��3j���O��B�C�GG|jh�4''�]��9���(�_�u׵�j������u@T
���Ryd��&R��5�wq�,����ZaOa�O���M��X�J�L�5�v�V��-��V �i��ei����Jb��>g��5���:m?�}ü
�Ctl�AgZ�?�
�z������d�v�ZN��y�=��^����1:�O��-6{���RJ���O���1�ځ��^h�]yI��w���p`s��7�����F �ӛu������$'GgB��ہ�;�p1�����c���V�j��qӊf`���E�4�%�#����r�+�Y'�
{����$i���{m��R�R�4�Ti��iBcͷ�oJ��E��khĝtm�&=��{���xg��(�b\N���k>y4�i�l���f:ye/�U����Xa���/��B�-beW�!��RP�-C]2c#dx�V�!�ފ1qx		n��m�\�LJ^�c!�#b?�WE�${9��#n��T��K�J$0p�o�'kT��ݵ46��cy�X��a%c�T!���FЃD_eM�tp˩�N+7����~�;Q��ܵ�%p���'�:����S ��<��Q��瘛��6�����K��E&�!lC�� _���t�����m���R~V����9��r� y� |�}�S�E=3z����.���$����u8�mt�DL!٢�Z�G!މ�S���m�`����5Q�E�aښ,:����F�Q|�H�}�Â�o�g��|��cJ���D�-[�i# �ݥ�R<����HXh%K{�%�>�)�3�l}����/���ҼQ��%Я:3�%b@��V�����u��s:�ȗ�3F���Iv��V>�}Ißό����k%:f���=�V��=�Y���"�2�(=L�驅cs�k!?;��F��:�?�хBL��J�Ԉ
��:[L�¾�G�"c�c��t1Шπ��)5|�����S�NQ�)���Q��Eg������rgd,L��g�;]o�}Nᥭ|J���x��m?P���5����poeٽ���d�č֠D^�%�`�nm���H4ߏ	 f+d�Un~ݩZoW���.7��kԌ^�
:�n��}�H���!��7�pn्cG��L�$�-&����
�g�j�r�m�6#��s�V⑻=e5>^�#���@��o����p����e�ۀ��,������tT��!��Tp��tq� #nĜT��,��r�U�1.B�43�R`�����p8~
޳ �F�#���g��b�:#J����Z�������!����A�%�1�N���gZ�l�F@M�.e
�����A_&ա,�=�Ш�N+3�C�ad��x����I4�e��^��m���Ql�pZm��ͥ`�jf�W��^SIW �o��V�:W����Ēs�2w)���}B�LIH�]�
)l=b�C�7��Dڟ��f�t��v���������;���I?FD��Ik�&�K�[v6��ŚO��%ˤڄ��1ہ��c� ����q3xS�qP��rx�͡�=n�%M�d����F�҈��݌./�4�x��5�A�N�E�sFA�4��~���-�X�=3���@-.��?� ��i�'����*�l���4��km�K�V<�q���oU�6;gG�H��Ҽ�s3�����		9w�{Ot(�*N@�NQ�t�,^��@�Mt�o�茳Oi��v��ڵ��K�������R�dq�u�Y��*��E?e���;d&�SMP�R،D��90�=��#�%��x�����wf���P�	-卢 ~뤼�й8��GŃ��_�#kmCߢ;�j�����{��Ε��d#�~���R�m!j�lwP0l���`�7��5�e��t���a8+����p��WvU�xF����4��!���h�T�UF3~s �Q���4 ��_�ifv�y�z/�u�����g9���4R�	��{gA����}_�]�kA{���N^�O'U�ת��NY�G��U�|��Y�ڥ w��(����%�t{$����l�n��!�O깒eJ�*ʰ��K-�L���<tK�恒/W^E��Q-'����ռd�`�q�����ʝ�k�* �JU�v8/�8"j�k$�fc��X�%BO�c���>l�9L�?4�C���8�GwIK�Q���셦J�W�zL�ఴ{֋�Y�S]}���� +�'�:_ZDC� �!w)�	s5��P�#`�e}a�`7]�����F\��|�q5�qp�nh
Y
i����g8��#��^<�[1��z+b�k���F0*X��J����C�����]r4�3�P�X�]	>G�qt��?��n�5^}��������;�(����PL�J�Fp�������e>�
���5c��Q�.EȔXui��c���3 ^����; � ����z�nOj�������0���=f1�k υ�w�v��K�X~����C�;���"�_/��t�vp��qҧ���?��
R��HW1
�+4���ۙ�!��b�����}��]9L��m�]蒁��̟Cr�<��y���/g��g��[\̟��b�J	jO!����!8�9A�W��ir���5~s�2��j0�ő�����Q}"O���V֯_Q��#��Qc������ek?�~��'ͣ�[r�)��S�����<x��� 'ڶ�Gu9�ǋ|������"c@C֮Q��C��j���.���]��) �נr�R�5�J��O��U6�"��cn��2���q�.��Z혿�>�[>ciYT���Hۍ�=ȩː�a��8X�:��a�w�>��_7Ύ{Ĝ6y(z�#Tv-�%��a��S��jS,�;x����K1n����d{Y`�y�c�#@���_���ҫ��
ʤ"h�5��ekm��L=�%#�](k�I�_�� ��Џe������n�ג��j��<����8���/�q[��e�Ղ�uw?JD��O����"G�@�e?��{�i�᯵p�"��dqAc���+���}��ô���s���[ڃn�����Z%�ܬ����g�1�8y�#�v{�3&����/�#�^��>��������x���{偹wH2���A����D�/��T��"	�eD���.�{	5�E:��=�ZF%��T��S�?�]/.��?���EV���A+��M��&��R�
��v�8��::��#z���V�$k,����TLZU�  H��8���龻2���o!�o"w����Xb2�A9I��=W-��W�2V��&��WJoU�e�w)���?3b͹@�(H�L��D=`��������8:�֐`��tdC���� o'=c6�\��T�#	��"D��z^Uy�s���)��B=�l]��X@��Mt���Z��bڶ�rU=��%7[5�M�6�̙Ō6%���o�9���C��R2"⅖���u���=��碸�v�0��ƺ�!�#����Eq����Gxܔ�Vn��#\������>��wxi����u�Pl�:}�0�Rg� `����x$�X䅤�pt��q�ež4}X�?3���^�f���
��u
#�)�|R��@I� ��t� ��q��ZVB]ר�e��KS��b�0���\n��y�5�wY�1��;����?�����zS�=_+&AE\Z�v�;t/9E�Uǿ���vE��i�-��c:ɂ����-��H�NW��A��h6�ol�
v� ������n1�Z3���ep� |+r���lQ"��?ʟ���8��Ó��}4#��C���3�I�����KAD>}����8)�ʎ?Q���q�lsa���(�<^�K�ר����:~!S��P�0�Y�mT��%��������2�z +>P���&���X��M^H�<��[�x�)~55�vE�?�Z߼rH�6��V}�9� Q�F� 5�(K��m��e*���T2<�����>�\�{Vh���![­`
�_�!�t1�^�>��
Y�����3�)Trh�U��5b;1��]�d�F>���_�reg�9�J'*V�$��`�X�³�C���m�U)�s)���K>}�%��EB}v�� ��uc�@O�[頧#����}�g:h=тLȲ߷����@^Ƒ0R�a��G��uh2y��<��	"˗�"y+�9��<����C�B\�L�uDf<e��7����8���c�h�#�]n[�#U$!-��{�8�����os�[G��=䤔�<��A��,.]s0��>#�˩�*��_H�Fʮ�+�E�;�M�wy���T���Y)�p������$���Y�I�W��w��0����/��<�Km���u�d"�-�)k�V� �7]�m������Y�7����!�����TYG��� �fO��n��I"�09��P��\	�TT���<E�i���͸M�x_Y�G��*{E�w�t�kÖj�z�
�f��0o���'с��m�r=��(���	0�_���T���	*��kh�J����x)���p���� ;����E 
�?E~+�>ٔ9�M�,h��$�Q���9܈s!�dz""��-���h�If5�n7Ն��rRA���}j]���A�j���n��?��UC��x�WD����6qM!���J˹ ,�y6��1=y��xˉx�ɬ���	h����;h�fHC���.����K_���*E�����UL�m�t�Z��O�C���]����k0`M�>�����Ǳxi2�d��J\������$��,9{��җ����1:ى��?�ǵ�нM�ʚ��-�d'�:�G�D�rY��?�� ���bKSϧ�\�mːv<��O⩛������\eSǓ�0�ʈ�5<G�'�/4���Ō7Dxd��@���E\�4���&.�΀Kܷ�
��s��j�v�}�����L�$�5�.:^L�[?�g$G�),�V��D�a�C��Nu��%,�H���(�KB�x����F�RE}О�?�1�f�"{��8}����Y��G��S�si�ƯH	_Hqm��<���o��ׂ'��attLN�덈���G�.fǬ�S�%1�˖���PA���M �!�_-�P���E���kji�	��Q�PU�|���:�e�ۆ�b��f�5\�h(��Seh�j��}IdU>����-ٰ#O��:w]�,�L*�)5�em��k�k	�D��Q
��1G��l?���&�Ե����H5���������+/�\��7@5�c�O���c�wv�+��v�`j��ǭ�{�-��7ފۘ�-�ج=���u������U@��k��<��8�Q˶b�s'Hu��r��6���p�S	�R�!Z��g�ttߓ���5�vO8��"V��B�2JhH+i�S��7V��<6U,T=�f��<<�'�I]D�P䎞@�@L�*{I�!�r$v����X#9Yz���o% �` �$�
f)	�{֦�ϰ.��x\��BC�^1{}�����!���ݤ�;� #�~^��I�S�������s�'����h�A\>���`7V�~lb<�� *���(UЧ�`��#���Ŀl%a��KR*��n���o�����C�?&�K�����aQ�,���b�L$��R��*���p��[X�r��B'����"��~�Fԉȝs�v۩18�*=_�����B4Q�~	�X��I�b�ϥ����Z�e|(
��|���,��%��/��7��Ѡ�7P���d���\:�Bf��;��՘2/�5m�����{X?Yn���)�"YMBF�ǗF��>,2iw���� (�`�O�@�Y$�V�@�H������͵ݝ��q�<�c�y�+N�q�~�]ɸ���y�g/�c�����m�%�L��5��0�F%?Q�OX�й=x���8��!��y�<#c�t�{�y��r���d#�0, 6�6�K�~Z��O�-ؠ}c�7�2��T��@zo��0bh�7��M|ޕf�gLi��~⪚�7�'S�ϡٰ\,[va��=W8%�2�Io��Qo��+w��I�$����޼�K���L���)u�5��s]�O�<��0���	���`I�b�ܦ5�1- ]d"�a����Ac��w���r�ў�����bhk�h�r���1(C�:
���L"3�:�O3S��n͖V�Ft���1e*�X�	�/�L�u�Wq�U���q�,�<Uv�r�P5o}agUV�{Km�9�藵��6Uk�̦� �����.��!'i�O�
SCEq;��Sov;Æ8�̖j��X1��Ы���z�p�o4b��Q3��~�
~]�Y��r�
ڏ�S�T�����4�8|%oi	�+�#�ˉH�M��hm��B?f�_!��f���y{�Lw� 9JX�B&)=��,-��d�6��]��#(��8�h�H *������[Y�h 9�����pM
��ߘ��5�y�����J~ya��*	�x���{)�j�s�o���NoRa���S�%����'*�},����7t�=V��ޞP��<+�w��]d+�3mo3nOP���- �OۦUu���y�F�Ǡv�/�#���S��C�JX��c���?$b	�Vc�X���q	|E�Q�9*;>�ճ�����zkR��+��m��"-ڵH��Q-�V�d��N�o�ͫ�T>C��0�S�R�����숹&��H��'��]�S�*y�������������F��MC��k;�N*lY����kC�M�; ^���d��M����r��10�d-ޙK��U꺫�ey���N� ����JD��5�%bCG�����5B�3>C	M@M�ߔ�߂�{F$�Ԗ���+k�Z���1�6�b����W�;�$b�a�ʣ"�6��㤇��]��$W��Q5�y���[{Q�(�Z�~���5�f玸�i����"��
s�~��f#qe#ug�����y����-�,��kN1�ԗgp㭞�ˤ}�N$Mq�N9��ɺL�۞��O���-%��L�Q׀��1��T�KA�E�������a�W����}G)H� R�L�
0�א���*��/ǟ��Զc�h5��[�"T+Kh�#���T��R��PC�4��(��զ���i�%uc���Gz.�#�>hB.�3�=�;�޺���bB,�D��q��rx���_�SHZ�r} K�s���M�<T/�X,Dy*�94Dl�Lj����y������Vz�T��6��v��wW�]?�St~>�?3L�c��9B��?L��6��������9
���C�)>�F�U�6QE���8#�b��=�����Y���=A��
���E'k�tA�9׺;+k���1U��M����.6\U��$&�f�ه���f�:dƒ.'�ZK���?~�/Z��A��^�I,V�9��C�6���!�f�'�$�P^�G>^<4��^����z/odL��1���vD��+������S�@��-���:�Pr�<��/���s�Ʒ�s��!b�`����#�W@���jVK�oUS��{<+5\�Y���t��	��i�-a��KT�d���t��n3[M:�*9��X.��#�,|���X���*J�0�V�q?Ev'f)M�I�%�����ܲn��#�J�Ι�%�>aTg�G5�W�AyéЕ��G�9|w��tzC�u�Q��}��*a�L5�]�+*(e�lE2���X�`��>�Z��ذ쵝��t��0�Iv��C�%62GT��hX�VЮ�_�u�Vd�ŤÕ����
��E���z��e,$q`g��m`�`�ke�U}\A�2����O֌�h�8�&��.tmW,�K�:�\L�:�"�5�ɿh�nb���Z��]&;�H�jEI���Ռ1hB�㞉����������-�N9�R�6H� r�$�?�, L��4�x��ث�e�IU6[ �.gN�-����ܑ�	�FyJ����`��EMp������PW%����H��H�yݱ���c?���o?���7�5�h�x��ק�O���zx�#�R5x��p"$@���5[�=z�+%���Bz�~.��:ܝ0�$v��Dan��8��L���]U�pg� %�ן'���,�v;� _v�s~ɼXi�W��y�C:���?�W��Ȯ�VEY����O�ܛ{&Oh�����E�&�>gC�<�_9� ����������s/���yB^ R���.R�y0{׆�� M1^a�U�L22��t)L񃴕���������3 ��� ��"��و��->�'ʏ����h��G�n륻GT),����v91oθ�W�X2��ڐ�beڤ��p�����~U���9HR��4��T���y�(��YI��$��#'��[��3�?�<�v���5!w\����a����ɾ��:�ށ��#r}Z_EeJ$���g����'���.�=,�������8�e���F��ˈ�?��H���5�5Ƒ�{$�����k]��ւ8iN��m ���UQ⭮�Ϥ����Գ�yȔ7��Ī"���lB�=�u8`�C?���o�ؖY�#�G��m*�v��e�-�31ǩ	��Zk!�%�߉�0G����3*�g�Z�g���w*�-�����x^rW]t��(�0����e�����*��7�t�~�-���F�~ߦiBUǣ`4g��B�	`L�Y%�{>�ƆlQ�N4�p�G��|�o�"��N�aOml��`�4w���n��Pte,���O���cq�W�	���wQ��`�U_=�>t�B>���n�n��8��U�WG�;�&��9?-(��AB�MN[_j������.��n���ŭ�v�lb�Y�����,�(A�@}Pt�����T=��hxH�Kњ�i2S!lQ=��1a����a&^6䢿#��w��%$x3�F��Z% ^g`��4���[��NIp�b�Лq!��#A�"�C�����ۥ,�R&�\w�$�_��w`q�]1��]�#�#��Z�S��ސ�[/�N�c�(��I��ڥj�� Q��x��I
�U�y}��Z��
0��eTa�)���8`�����f�*���	���@up#�x������N�@�7i�T����i�6�(���Ӷ�^Ժ\-�U$���~3Ԟ* ��p���%�Uiq��|��z1�hw�m�=���KN��qr��I�n� ��F|��xE�9��B�N�֖H�>\N��uD�%�on[@������5�1�/'���Qu���'!��?.��
��,�@�C1P㝓G_�X�)�3ǎmh���� ~��;����F�q���Rm�8	�w.~fd�q�[� q`��-T:��r�c2�a]����7���a�#�b�U��O��M~ZT��ћ:s�	ߧdi)af�y��ťE$.�C6P32	Щ��7�D�o��U^g��8�T��{�$%4^�+֋Y��e�b�o�+�^��Y���5�L���2��p�z����<u���aa~�$��`o�p�#��L^�\��s�֦�J�ϳ�yr@P�}g��]���ï��?���z�J�� �=HY�.E��'[Eu�˶#�OR���ɝ��'�X���[��!7��9$�f8����^O�ʇ� ��^��}�і޿�n�iɋ~�<W�R"�k>Gs� ��W�۶��m������w�픍{��r�V@#�M�T�Ϡe�fo����8"���$I#AQ�x�p�;4���Xu�,tS�� 7��x��`Y�ߚ�oq`��N�|������M�1�g�H���B�ǋ�"P�e��o�r�#���ʹ�b���i�H@5�H����+6� o����ߠa�_�[A�a�O/d����Yp�4c���fH �ءw�s�SÛ�p�)�j��x���1�u��K�!��F���.XgzX!���酂+w���F��bh�x9���_�2@js"y��C:4Q��c�E��!E-z��W����I�!-���X�t@�ϼT��G!ء�B)�T�?�D��H�ٰ����̢�S������M����TQ٦�~���j�_��?�4+Q�'A�V�உ	>-�I��V�?��Okbq�Z8�Vo�ظ�5����N���7���lb��7��)�W��{��C#�q�,��O)��sO�+�Sm/�k'�$�V���3�XBc�GK��1�ñ��>�T���*��I❞��r��5�C�g��)x�ܦ�e>�=w]�=�w�� ס�m�9��cLM���x|�P��٣m�f�2mC�ڤ'Dw㒵GD�6������Y�N&hvU7<)��m�D��N���;��E��}���o�L�[�L��V�<��9;yx}�?��0Q�7�E�F�)�U(k�Zd�'ޞ��q�r���N�n���1yAyKx�ٗ3�3�Z�I�O��4��e
�e�E�SOR;]�y�$��,�5T�sG����ғ��v� ��^�u����e>B���3��$�}"M��@K����#��MF`q���R��_k�D�����=�O�,����A]����ĸM�*����p�:oդ��фήP}y���J��WQ�v��o^U�o��6�[]���A���Ԕ�!͒����u3*�cgtܑ����}UD�A�5�:��1��C��A!]/�� �@\�����!�����aF"	
n�N�R��ޑ*�)��+p�k�N�gI�J3���6�hQ`z���f+��d�GW�1����,�W�Cq K��[wk�,�[:��r]}����G��ɓ��3��$}�z{]J�HO �F)I8��?3�l��ੌ�ۀt�%|?�7���Hx,qI,C�qfh簙��.B��&ODz����"'�cCg,�����R&xR�	����!0'u��Db
����fk�r$��o����0e��F��#��hęI����v�N���-�T����-~�ك��^�`i�y�5��f�<��5F������ ���N����ݢl�^�n\���z`H@<
br�[���՟Y�����v��]pq�Y96��K/�.v�X�k�����%@��p	a�ږ?�1�k�#�>�e8�"f�%O�+�V�+��GPi^X���i8�B�I8So?L,� r"�Q�*�4)���X�� ]����}��K��w�=i\���z�PpK�[��.)o%%�iex��u��g�V_�v�C�[��t#�i����.���A�R�>�?�%:+4Z�ߛr�L�V�i�,�:%���B����cXIk=-�чA��:j�'
�2-	�σ��8�����?W^{�����r�G��/�;�_��EN�f��6ٍ,�1ɞ��J^T���Q��l%�Ϝv.q�5��X��3j\ S���#���0�D
��1�7��!�y�����]��� p�q���p`�ġ�k����)h`'dX����&��̵�R��M���ׂ�E��*��d�y�_�P�~1)~C��!`/�[!�����lҙ�QɈpx�#� ,4\Q����jκ�Í��M��߻P��ʓ ��x
�8g��yb�{|j��W�M'�Q�C��RF���Z9Ӽg�*�` e�7�b�hJ�Z��3Q��T�g���>ɦl<U����d��o�Ă��_���ˤ�f�P�3����1v-�u+.@��e-��M�'˅:Y'����񮹱o� ����BYUu����n麜� ?���w ����R�@HQ\����y7S}��-

�%Kp/�2rey�b�>�;��~�Ti�����@Qf��j��[��4��f&�?a!{��뻧�M�4�	�˯8y1��׃����h�b����)M�ܘ5�tn�ŕ<�FB�q�$��Դ�R�C���FڢK��u'��QQ������9 a���Yd�l}���v����]�x2�M���-g�<�]��0;A�
�/�kgս��c���?��QǉyaX߫���L���eO�w���E�v�J���������M��/� �a�54+�j{��؋�	t�:w�y���`U�(	���n�J��?�}��]��s3	��0:��ұ�P��<�����|źa�`@�G��PC���o-���ٿ4$�/u��eM���&�8T�o_�P`JNl����(a��&��Z�*�Я��S�DT]6���\#6�:4eQ.a���v�R�;{(�ry��).dZχa0������ �\�8f?ψ+,�s�Nm���9���}���~@��"Ҟ2!֨>���O�LW������,�_*�۵/��6v�%����ܻ�R+�0���<���?������8_)2�+�@��?����Q�b��H rjު�H>}I�K}k�;I��e���y͂��$�e.f._��V�̼��0���x��XCQ�4�a��|�ꕂ���9
���5��g��e
 ز���LbD莞&1���d���3a�4+�~G�KE�V�!zM�H�2�{�p�/�����+�dN��i����b�v�I���ӫ�ɜYu��#��jf�pZ����H��*���HCh��hwo$�#�ǐ���y���Ѳ�y����ڹo����U�F��ͪ1�8za<�)�d��҅-�Y�.&��e��K��t�g%��d�َ\��;�J��;�s'����1�=�����I%J#���� �J�~��1w(��٩0�x�Q4(�0������6��{��6�|�"�}�ā�=�F�3�t�-���I�B)P����\
M��a��zx�9gp�9�E��-ƞ@��<)��&�b�eN�âю��~"��������Ph��M�P�^���$��@�O�8]_ql��&�����ń��,��L=�`��~�b-/aЖV���k0����n'�a��r�L��ÑH��j\2�1-��Z�oS�̈����iB>V@�Q2�7�WA��}m������оY 3>�,0K�4-I���9M�QJr�t��������uJbf����^�n}p��s\����lOK'�A<���t�a��5�x^k'k4�3�ց~�I%gСs��/���H�e��\{S��pw	m�P��bńd�W�I[� ��l������u�=����,�(J:��^�`pdJ=�TwF�d�fz�`a�����_������F�M4n�piP�`k�00�8듰�@����/l�-/��&�4�t�z����Y3���č>6���V<�^<��ki��ݻF�%|g��'�i�p��U��-P�и5��^!	ނH{��?`Q)��1?����P��쾂P7F*����{3�PBCC�_c����9qN�db��u�~
����
C'�xB�������ݒ�#	pϗ��۠�G��<�=�GiVK���C_��h�0V�F	e&'JX��J��_��Z ?쐌ʭ��YI[,:S��1����OC���5��	�r(����6FX����xk��G������2����@ P?'��� o�lV$�_�E�҆�w�.eCî�Ĥ�|�+����b4i]2$'�[�)ⶸ�J����w��n#%f$�t�Ԝ":���h��*��޴�<�X ��tt()�*��2Rr��ʹ��@�׸>0d����I>J7��������_P|p
�n߾d� fv�e>����7�;��6}���OY�g��6���$8��R�&�f���"Ԯ�D!+|n�����w&����hH$G�x���ŋ78�}�t�������`h;7���x[p��s?�]�b��-���>��ggَ,\���7�t"v��"`�^�Tғ	;�B�f�y砱H�]!x_�!� MD��e�*�@�����2��$$�&�U�{X���c,��j	�"�Ir�K{ �;Q�,�ܑ�k8�¬^q���U�"%�[k�B]^�vg_bh���� �FvC�r#�xa�y�F��vG�p";W����[ª�	����D��6!�� ����E���d�"]r�^����YE��g��ʼ��g�f�����P·I��k��~���]��DY;��u$�(������ᾞa�lL������o5Sa>��'2<sV��W��h�����#�Ԃ��/�\����8Y�
���0�qK�|��ޫ������1{�=n"�*��V�#_�]7]+ܗx`�B^�[�@�+Y 2&^��G7�q#f�_�G���C)D����I��:S� n������@�m���G�m�=�2��efǸ�:��uK[g�B�B/2,���6�b�~�~�����X#e�o�N�	�vRH�T�R�4HD��=t9�_n��1	ʶ eCC��0=ʺI���Mٚ�ѵ����,��i�����ʹ(���J���һ~;�m���5���gD��C��O�Hf���Hq��,�;eӈ]#] S��<�oMd\^�$j�L&����a=��.�p�̳�8�X�=��M93�X��zZ)cQ"~����)�+�ǫ��"�=+�>�9�	T�`i�l �(#��Q�z��ś]6-H)ې�S�f��i���(^�7"����毡]���
�-n|����EҾ��|�E�M���ډcֹ��m�1�	���bv-�l�tSYgd��!Nw��ϋd! �������:\B�nm����ʊ��i�S�V
��R8W�ˡ.�����IJ����ph�M�%��a��if�޸�4����0�q'>u(R�N�z,Xg��az�;����v�Zp]%z��V���6��aﳅ8r�X�	V�[�������8���+�A#��
���|�-���,���x�\�Qok.8�V�,,Hh+cS��%���v�i2S5�*jj;��h��1�E|�?�m����n(��&j���Pn}.t�M�U�0�rf+�vB�>Wj�C;�k#�y��B%��_��e�����z��mKG�E�2d��;Z�b=�k���*Po^T��l���w�{!&�3皖�
��;�rqW8o�4��Ċ>�\H�?��V�F#�B^=<)�o�q�s;�R��'R�r�N���_,�)Xu
؈� �ϱAg�&M��0]z �xX�*Xc�o�8��'�E�����O�EP��wk���`'�y�̶��!�����$�*�qx��o�ؔ%I0ڔCUΰ���n�f��	��9}Uy���T�G:X�1.���VM]�mUa�+G�dL�5[�0��d���Bi�Lj��(S�oM4.J�}WA:b�0�c���#ˀN&�`���T��㽽��{	�]S���官a��*ǣ!0�>�lz3���u5\!�l�G�˾$�y��
�*���{=������wƂ?�Dy
g/"��k��:�t�3��S٤�E3q
-?�7��\ì�'�yj�w}A�2�O����}ژ\&��et�W��<N�	��B*�]��0�iC�J9?Q���`�\qQ�'�5��^,�p�S�V=�v�|ɡU��.�^`VY���>AJ����mp��C��K�k/��&����&`�f��Ҭ�0�x��fUo�mB3繹,����3`chHp�Ɂ`U��/��SS�67TwBy�"���t*+�v�@`�����%�����X����8��3�O���8�����'��-}j�NoC��Ӣ���.p�u�9z�{!^�k����g���O���3,�oo#n]Y�w��zo$p�bt�vmC�g�1��*[3K���5)�n'��%@�nw���1T���]�\�Wef=ǋYS�Y�oO-�E녌@�����Vб�)h��n{��]� >�D�\Ǉn�2��@5۫1������Pwg�vt���D!B��Խ�e�ea�=Yl��Z���u�;n�b��F����.%,-`�T���w��l�:q����Ġ�Ȫ\��e�o�H�7ȥ^�3�"KV��������B���(x��P%�1��]Xr�<�֢����{���GM�c�A��0�O`yE�"d˷%G����re�ʠ����*&^�U��L]5�E�i��?Gj�7ų�_$�f
��
�B��o�6eU��6�j��#[�!Z�Yv�A4���Ly�8�����zn[���kf�r�Py>_~Z7Ј\����m Ê�9i3D�nN���8>��&V׶��sF����#�#AQ�M\�%�T�$s0Zų��8���f&�aFg���F�p33z�/�bn	��M p��l�oa�/h�"�zb�����6*�����(�K��avM��OYѬ�d_������~)91k�@�2X��q�1sʼ"#G�/�}F��p���� ��i�*�;G �[y����,v�2ɻ�F�V�����dSƃy�b�7X&5TM�Bp1��3����RV�� :(��_�-QˠIY�fo��o��#���C	�`ś��2������r���=]#L<��m�E���Kq�s�$�Ig"��Uft�ر�I�]�M:[âǘ�7�<TR����Bh5���I_/�
�PUA���S���{��X_���0�u�\������T¦�m���O��aT�+K4����0h�yĔJqJ��` ��;�Z�����Dz��2�Ģ��UơJ8�PKW���>J���?�q�f�",I�Lޫ3�	�	��?DߕǍߥ�jq�n{�Ve2���6&@�4]�hx��>c���1.�����эY�U���yx����QvY���f@>eOlA\w�v���rA�U�����F��=m�&yV!�z}�{*A������������v��EÉ7) ��+�({Q��œ|��(Q�!��ٓ-�kW�`}��3@q⸎?�y�"_H[V�sL��WDu���]9B\<��a��[�{Q�V�)CZP:�9��"��k��^C�TjL�Ie��R�3J�q���ņ�/|�sZ^��`@�d�l�����>���<��gxُ 2�@w�gmD��E�$Κ%9�V@naV�\\m:ˑ�����CwfC�#�[	��f�*�	F2���)���;�%�u��ר���B>�w)A���m�1�Ś � ��r'��re�"Vʃ-����C�P 1�C-��V�y:�GY2�|�?���sY��s�Bs�_����& J���~�R2P5@�[%���*�z�g�vȯ� -vE���K���C����=MA�gD�"Xg�[�F�r���<�����P��- �гT>m��7�'�v���-�-v�.�R)F^8��h�O�'de��q�Q���t�+o�Gu�G�� �G��n�+녺�Uܽ��aEm�g�j��^��>�������m3��b?D�s�w��������գS�)2a�gb�3�cs�7���pp�GD�`&nGE؈F� j�d@�H����� �]�J&'r��Rw���rH����5�\��ʄ�P�P�v�A�!膁���v��� w��H��\���j��x9,2J%���`/��,�z���lv�[i�!�PcK�G���'	���&�7Ta*�2��к!�W�����RBrL3����J��@��Un5��p���*PTl����@I��cCA��es�"u�p�:�Y������!K�Az�G�TkY�ׇ�[wF�,��s��\�^���4͚�%�#�L�5��q�%�\^&T�U*�+Q�>�Ϥ��-�JFf*g�'<ѽ�