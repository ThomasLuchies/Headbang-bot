��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k����W�z�N��VXi^�p���d����So����SҼ>��>?P	㞸a]��s���$�Z��a�	FG����fK�n~��|��v�������5���� k�ɤ�&��d��7��o�$�,EV����I��z��$�gQ���R�\p��\�.��s��<��ԁ���rs  :���j(<
J}��^�U���<OѴl�bŋ��f����Jq����C�y[��Sk��h����XZGI�tU��j��?��J�������	�Nx72�n���Є�(��슅�V=�X�P3͚�S8&o7.�nX�h'M�\�x��c_�k2��s�����x"Ux�2-u��hE���;�(�/D	_�m����6xD��,
RLZ�G��n�"�ݴ��Oٶ�J8H�����O�ޝ�'����j"��D_@��q`Y�SDxgc�a���>��0f#(O�?��
��ű�U7��+l�-Y�GX�u�eu�<���,���R��ꏠ׸�龠Vm�v�Xw��xe�A̳R�5��!����z>����9"(�|H":쑊��b���b��w�������:�1�	*"����oߏZ��׶8��?'��'�-��Rh�ǿ� ��H��#��:��$LJw����H[T�U�Ӭ�j���EI��+i�r���#���CH��$�a��Y�= �����7f(�-%����q�A���͸p��+�\���&#�HM�ω�NDV%�]��Yl1g��k��{;0 h�ø��!+�˧����4ޢQ�¿�;��-�(�pa�y/c����'�0��Dp�����f@�c)������c9�;��*���VVhVc�U��DCc|�\:[�}�	�X��������# Yjv,�Z��K���{�;��
S�|����\9k_��kc �h��_y���F&v(o��6ˋDn��5V7�	� ao"���i�n�ۏ�: z�wO.����^����r�S?jq����������Av�5�FڻƼ��� qVx���6�|,���Uۯ��>���T�vM�ŇO��#���7���Q߲��ܸĝ��+��amz�1�vx�jٿ!f�P`��Ӻ��v��2F�x��<�����T�'�gqI/<�*�P0����5Zv��:�w�wUHNa��vP��=X�QP����Z��R��q�Y�8�@6�I
æ�1����m���8�{9�y����rǔ�!�xa-�>7�lOlХ�?!4)GmZ(*`cl8����(VO;��I�B{ϱ�Ç�P��3t����cɶ��M��g.۲�cQZ����p=�>57TS��G{�3g5|A���ub�X�z�L��Sf�� ����'њ�[�Ո,.4�I�w}=�'(��\���(��I�:��X95pLSh	�~^X�X�u5��`�	wN��r՛��^|��Q�w��ε��<�}D�
�L�F�>�>��o'-]��tl7'M��g �@2�oב%�x�౗�R�a@�k?�	��B�w�̬���9�3�>ٹ�a����ײ�^s� d��I�)��rl�F(@XHV2��F0�Cp>�{�s�&@<�{Ha� ��HئĿ�g�|��WJ1�|j�_�u�Y/�P�[z��	Mtn�mx�2�85�9B ��ug� ��;������G�����|P��j��aL�)<�B�;\��0�G��vOJZ����Z�.�݀��p�(x��rW��yܼY�lkLMM����Ю�Rw=gS��o����㎏�<*k������B�x���� ��[��I5{F��-C�2РV��Vj�w ��\�ۛ���L���s����7y=�^'��D�;n�ڇ�bhp�&��y_
�y�� �q��և[BBX��G������P )n`�p)��r�\$�q�Yo����p�2�Tz2o��J�}���n���	�?1=b��4��bpd[t0��Y��	��G����gk�V2'�k���q���^�5�^�^�'2���/�c������ק�&��^�d!�Q����i.*���ƈ��)�yfUO��M��sEI>Q�@���:խ.���tϷ*[�Q?pY����f$j�@�l�:,M��G~Y�N��uѵ 9�!2ؐy���l�r�.�� \�J��[��,%��(7����=��a�%����K��@��Q=���![�}��'�b��c(3���ߍ�?	rR ��n�4}|�7R � e����������Ifܲ-�~#09}!���n���s4X"��~y���Z3f�0݄�6H5�RW�x���8�Y��Έ!79}8q�'7|�B�����S"��eH�6�����!�����'ފ�ʨn̗�����-�~8�2|H�H;����&eS�~�M�p�7L��`ߍ�,/,5kG�"��T8I�:`��6e�X�V�B&U��h/�B�<��v~5�%񎉥���%X�V�X���8<{˂�i�;+U>[�����@D���Bg�S�x4�&Oė�t��$�0E�z���]�|#���՝�LDţJ
�d�lj����!�r�>+ɟ����$��B}�i
 �F�	п??���tuA�?��eV��qzߤ�u���J�^Il�i����|!��f$p)�F˘��0�n�����6�5]�K�_<:�P�ݠ��:r!�����=��-ן�"�ؙ���T���Y ����WU��Xܛ�����5Jq4�O�����������?�RJ!�ďS�b�i�?�����1�w�h� ��rf(�R���^�Z�k�$SۼLw�67[f�;l���l�}��CI�Y�O��
ߴ)�q"J�Ň��	<�,*�ν��1�W�F	��l�����}�駴JK�ٕ�KxUc�����n�F��]���763��k�Z�i=a;�5�OJ�c���W;l���.<�2p�}(�n�tq�\�=(ڋ�$3'U��>$��Y.*ְ�$��+�&x��C��q(z�ѝN⭱�޴N��s�Z�i�)��������nTX`)��x�O�&ny�y�!���LBz!h6��D	(N ��wf׽���t�$�f�[�7�y+����#{q�N�[�TI�8$�,iM<m���2���ÑL^�)��ooB|�ߐG	Щ�U-XO�]{�4����f���AM�pw�F���(���XG�$ۛ�bMb�b>�5�:T�������<�9�JV����8�� a�z�PWnl;\ܭ�(f$'ӿ �p��=7c��ٸ����@��V���\�e<�_�їÍ:6CE���CѸ,^vC>>��)Fp7�4R�Έp��7���vf��D�`/^�Uk��:N)CR��Pj��ai0z���f�|��%MEg��t1вL�˫b���^�|��56����H��������j�u1z��pM���*Ŕ�Qʈ�F)���X�X���(�_$Ni�r��;ی�x_��,8Z�;B������DΛ����舢c������.�k*\��m�r;V�H;{�^��n~��
ڕ۳�[��%����ĵ����+��[���NT�� ������!�-�0y����)�0;~�r�R{j���gYmV��e�x���В5N"Ck�$�qى#8A�C6臠 }�mPZC;�x�C.�%�G����'�2��T!��� B=H¢8k`���
!�W=6<�]�����+G�X����H0L_ǻ�#*&C����T� �iLi�
r8;߿�f�P���l��ՎN�u�4i鎤�;�oHohpq�:~0��$ٽ��3�=�i����Q�4���ħ�|/��z)��yD1yY�Ǚ$�� |@^���^N:NU�2Zhz�hF�9�-̥�6?��������c��u��O����}�V퇕/�Q����>���hs�z[��A~��Ư��I�V1\2	<=x��aAi;؎����^����x,��	=�?H@��P��C��r.��6��Ws��ϧ�M|ɋ	�_-�i&�����o��Q'��U����{�-W��IS���H�G/U��-��U����Cx�/��Dy���Q�5�&��tNjv��!����I��U}��sG@�?cиc�n��[���7���F+�8n4��ʴ��I���#-�%���b'��J y�M[gb/FE��������6I�ҵ��Y��3|���`30	%E��W�Ʃۙ���ݶKRPxM����FWL����������hl����Q���ʶϫ�	��oRO;����(5YDYn�bg8ՌH!/�Bi�o��w�F
VFX"?�ž�S�H�������V�kY]`�l���W��4a3׫����u!(�O�F�����0�����y���=f	?>�K�?	ɞ�r4L!:"��٭�7���<4�U�yt=�!7`	����c�_���������Wmw�+$Ӗ5�cn��9��N�"8���N��	�����6O�mǛ.r������Jk�VbUmu�qOr�O@�]�����2����n�D��?/rd�`"��%_��F�J�f���@�!`J���K]N���R���`����4l5z���k<�����)���>�zt��U�
h]|� ]9lY�P��T��᭲�ʦ���1�q��_�r�Fd����lg�)z����,�LC��6ѹ��UuZL���M��N��l<B��faw�"��Iǌ��$9��C��͘�y�I۬�U���yH�ěk���&}z����ܓ(2>��DF"���A	�����r��q1D�m�yx�v^�k�|���)��\9���t����PJs5��Zw���-������_CM � W�?	��ѱq�5�r�
�Tn�C|��m�j(���K�D��v��9P�4m!
�#r�/�A�@`��Bb�CӓQ�v�,�k�p���pٚW	>�Nc��ܝ��F�z�r���H��>��G�n|]�Xq��9.�K Tx#-Qe��@o�P��_���n�����}e��;&u�s���oVZۄ��Ҕ��=>.6=�y~8���Izm#E���Uo��vO��T��a���G�=6��X~dTڧ�!K_�qR}Hǌ�s
T��	~&����j�	���ZE�!`�����(�Nl����Af	{����BH�D��Ÿ�����B���Z&���#eV^@�R�\�Fa?+ţ�U�d��u�;X���g�T�l揗 ����J�62��1��E(��E�i��PL���+���&�gU�%�-8 WZ����%����.Yt�A>-�Ir��1�W�0t��im��z^��&2t���n�o� ���8eMr�2d��xH��Bޛ�'��H���jׄ�	�8M�ط���v��5C*�mɘ-G���>�m����g.ԗ�dRޢ+�'zX��x����3�����5"���c�(ϑ&�
ǎ1~��VG$��壈N�TA:�R�B9��j���4��9 ��/�r�"lsЋlH���f�2���Ab�@$�\����ޡŏP�ۭw�8�Py����k�H��FyY�Gk����L�Չ�&fk'�D1���6�ܒ��N�c?Ը��!e}<��#���b<�h�o�
�����f���y����F�Z���[����7�QK�K�� G���+�h�8��"G��TǤɒ��e3~z)P����"�A�[�ݜw>P���_�q�K8�,��ȣ=�ϑ�J롞G��է$L��wg�?+I�)!�b5���OI��8�5�C�*c�m��Z*K/�ᑒ�u��k?a�Lw>�Z���#��ʕ�� 8b�POe���Q2�\\L�Z2G��́��ߏu�|�M#�� -	��qi���r��I{�q�q�=��{:�s.���<O��ߢ���L��3�Z���?A^\=�g���H����(��{���ah��z�2`�?<|Z	�i\�\sؠ�s��Q~�+P�|�â��= h���S�F�qN��+9C���'v�Z��Ĭq ���e��g��-3���Xk�ާ��?#}��Y���X���b��tt,?��$.�h���fW�����ɫ������s�*�oDY�����F��~��6Bz��źXk�kn�'����B:�O�.�3��2��/�� ez=��ZE��R�$��#�[��G��%���\�M+Lqz���6b�B3��o��vׂORgI7[$�������֙�������t�.��*M���Ѡ|����?Ϙ�9����8yL�z&]���'?�+�����9�GW�̚v��Z즬c{��W�l��*��~��Q�c핋�#D����d����	�<s� ��`�}Z�L�%�\H�H����%���7�6�Θ=P �K ]l[���mV��G�-�n�D���x$�K&�Kw�ǣ�	5�WQ���pHՊ�/��ȃ:���bK0 �a���ݟ�S�b���V��U�<�M穌�S� ���k�|�x�EOQ�I]�Y�Dd TL�tߺ�*;/�wi_�4���?!�$8;��r�Ɋ{�I��W~-�)dF �r�
sWQ^�J��ԳVHpO~��`��E�/�o֕���n�����=�������G�g,N�V5=�wͧ�B��2IX,�Q�O�^skًki%�_����l.qb������������ŭ�l�����+��"�Si�Jf�k���˶P����(�~�<��8���;���Bވ��IqH�Զ�4�V�\:�S�B��Q�gSC�R��w��PP�å�E�����t��.��(��#u\J�rz��f���͙W���ˇ;�����f�����}�a�]��2u*��R�.(�f����D�=us��uQ`s�[Zh8S�݂YJ����]�kU$?�(�4�|f(��k��^�������B/o�Л"�f�j�y�1�`��+l�݅��E���ܘ��s�xu\o4x�=�\$�Z��g��ȽBI1c��\�RXl)hA�	xk�ř>9���=� �>�����N�[b}b�����ds�s���$�-Bm�fG�֠>z�$�;9r&G>�52��s�:����X�^��Jf(Uk�%�B�{A2?�g�
�
��2o,�&xN7*���H� N(��� �A�Q���&z�������%�i[\��5��4���h9"�H��'�#΄�X�������Q��N�t�3e
$U,��0������&h� �٣����Y�sg�{_0������,/�G�Z��?i�g.�[.B����<{1ֹh�l���*+�6����6��;R�o\�-F~Ë�<�����,������3����[E��'�r�"M���p��{��࿺�[�;�V��7�pI����9�ڰA�rT�g����E�80aü
$�;���~�$�#�W��k쥶�1�/��9yd������ؠ��e��3�*�Z��hOg8�Px��ۖ�bB%l��U��g'
h���7�X��Wlh�m�'1�
�Ä97�j3Q(��k$2���e/f�AX4U�)���+�����9(�x���C�v����fS0�g����2f��u��V��k����k�A���T��%�;a����� H�}ƻm]�O+uqmMqsW�M�T͢�H�������|�wy#7�Q��,���u;�*�a�Ģ���'A�Ղx�ow�.|ү��v�j�S��!�q��W�ۙ�ͱr��2`���e��NzXg��'�V�v�GUAcU/>������u�x"��1�y.�E4�"6�OƧ�ۥ�]�fq��!f�k&OW[,�O�Æ��x1O7�N�I��z\�:�}�f���[̞TN�d	y�f���]F��-�V�T�d�6�_�4~�����n�uڪ�B��v9�&�0.��H `�dN�=t��̝e�E��<������D��`4��p,����F�K��q�W��d%1��m�T�����~1,�L�=B Oꬠ+�L�X����r/
�%-V�qN��~�-NT'Z�)����u0qMȦ�?�7ܱY��0(Lu�HO�&e�d�w�^��*�ez#�b�C��H��"'tڄ��6���Pu���0��c����-�n�N[ȱ�>�G�LU/4n��\6����{r{�&6�}PZ`����NxPE�� ���̀yow�e�k@m#��>(�����xz'?9��H���UWxP�E�g�(���P�/*9�ǁ��3��8䧤n�d¾j �# Pф�����c:�zԜ���\#%�	���`�����Tx�b�!�Kjɽν�d���dR�+��̈́`.g��
9MG64L���_H����F�،�Q���4���ľ���\�M8U�%��t�j�2b?oB�\KR��m#��?Ϲ���*���%�X7���u�K��Ϥ�������m�d�d/i�B.��3"{��8��ͻh�n>�5Pm����w�� ߭%jс\Nr$iRpDJL����J��l���'8����Ke_���Uxb|0����U��a�T��)pd�� �ؒ�ĉ@���J[� m�ג�d�閊ֽ��N�1�l�����I '��������Ey��z�.���$<|�a2�*��>�P�/���B�.Z��!��a����΋mmsιNޝ�U`\;��?�,`v$�,�`�l���)�^�eT�ER��[HH���3"ZzQv�[B�g���:ˡ�Z�����쉵*������aL"v���̠G��=�v٢��>���䋲��%i�l��ϙ�ѻ����\��`})��"�ˢLA�<7�,�L5^q�	
��D�%��^�})vb$53���Gez�/��L�
KR펕��j�1���i�B��N�T�w��&,2F����J�[�����Ǧ<�5�A��F����[s�r#G�o�Q�j���]t�g���׵!\Vԭ����!'JS�.�~�_{�k�O��+m�NM�KF��`��ҔyQrd��Q�D<p�d-֋�+'�1k�x<k*�>�Z#8�K���� �3�¿��UR���wR�`~0�թ,�3��V�/��������O�D�L��n�� \�'ʥ�KK?���O��50�J�C��U;L���`_�4�#;��`�v$��C�� ��cYt��f��UX���-��� ���!�����<mQ�heڕRVi�#��/WjBW�+�0�qN�	@q�#T^��,L�Ȅͦڕ(&�nGژ�.��m芄Х�p&	�xmB�Ѧ���5a�꾝��|/�������Ө	`�CV���J<l���C�o�h��賂B� g|�ጕ�)�ҶݑV"'�/�5�=_Q��$T���V��Z�kS.}G*�̞�����"�|x�_��i�d�cY��:#�O_��\mDۋhΙaN�0��D����|�;��o����R��ԿL�{��0E/Fx��`ʘH�/��gCI�i~BPe�oqG�%ie�
���6Vמ�7��vlһf���PJ>Xm� �����5zUS�+����U���:ͺ���E�D�S|I��������h�a�=�,x�,�b&�S1d,Q`o���qkz
Պ�V��2��D����q/��,�?�(�H�`^�|������NvI�~��:�� ���s�}1��3�z�NL����:��&�ĝ��Zd�*�@br�9�LtGX=���;�`D�6��q��:��V��a�s+l���b�%�-�?�Q�Q�>7�x�0��F�ʸ�g`�s$�v%������!X4H�d>��\`��y��|�����#��2�n��M�a 5�h�0G��� ��NGp�Cy�K7�\�Y:�MAq��r*ŊT�(q?��4�[�$���R��U��߶���\{�[�phL��J�H�;1p տ�!��qO�d~k���˛�vJ��ŊJ�K����)C�N�"ʰwrm�L)g�XQ�״
���*���$�i�&��d2�(�����O׮)�����FJ6RuWa�&�`u��'�g�)��j�>��H�+�����)I�Yʴ������w���ܐ.�Z��ڟX>5�5+owS�N�L�ǉ�c~9U,l�DJ�@�F}e_����HQ�R��"J=J_4�R�y�͡$�eO�N�7r�T�BŌ��c[�^�#�[(�[8��۶��Llx���Y�N[��$E���8<��������"��H��U���=�K�K'#�B�wN�7�L���E�M�G?{vo���2΀�|,j��$4<=��A'��l�Ѱd<X��������B+b� {��:s^V1�Q�.FP����H�k���������Q8�� �b����V��Dr�1�( �� ���!7���X������n6�-MZ�����p�k��+-�~B������l�A�s�[J���{h@�];�gH�ܡ>t!�y��w�Q$��f$_����s*�;���P�.�'%)�خ�lw��Iv��WLAE���#�>�̢�"��m�V;!�%=����u��[�E��Pn�)�RQ�~���.P�A��,�y��c�����J��}�s���z1�ԾiM��{J�Dq�
����zK9��3:;������"\p���.粍���W��� 0.��Ǉ)t�7��>{&)��R٨2!8�O��RM|i��B�D��V�n�{NE����[����ϗ4��;���ݸ�ʶ�&��*��$,p>INV�P��a�Gx-���]��BS�w��A�C��?�b~,5�Y�����$��~��8z���M��J��7�Mј�Ѝ:�<"�����.)1���`��FZ y ��Rg��]-D�����W�����c@��`��?#���b�_�ְ�簟��%]��`�d�9q�Sɑ�o�����\�F	f oZ0���.��;��r=^��̍0�I�:��ǹ��j����B�d�q�r�s��G|�����/��*��;��;� �X\)��Z�QT�7�VS����~,���zg�S4c"0��|(ׅ=�ޫ�xA��;-=�F��\L�t��Y