��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+�������;���ȹ�v{2� ۝ߎ#�W�ӂ����ݠ��>_g5���t͉□K2���Ec�ſ��`\_��cW��Y���NB��*�!�#-/�����0�����e	�.ZDG����g/G�lз������s�VS�]��	�_,��ܳЅ2꩙Ō��M=룯+�&HfUk�@��%��.���cm���pZ�^�&]C��l�QQ���UicM���*�qz��ZU�^u]�2�=>���J��מ�#�^Ķ���l�\*l^���F��A��N�QI�������T�xĞ��pǚ z���4��)�7�z�wcl9du�f,u���� OK���ي�H�I� ��l��.O � F�		�,& �����ͽ�`� 7�(������,\��S�!�4��ݮW���l@����1`q�f�>�U�g��E�����a�md������N���+���+���}���t�
I��-�&���I;c�C&�Q�J���5땕�?�Z|D�YP��e�|*���#܉B,��S�(����L���͙�p�&d�d�d;B�Hᨷ�ǻ��qa�+���  YEɃ��)=��������Hr߈�/G�S�>������`0&	�wu^+�#C)H�C��f�k��U�lv��v��״KOgC�Ѯx��X���8�xh��]�
�J\:�68i���Z�O	G���[s�B:�E�6M�x=	��Y�hw�946�֊0�緪&�td����q��)6�wqx��L53e�ș@h)�}Z
{�z;�L� �HW�o��>�������T��Ք�x���W��#�϶�s��B�t~��%B8��S�96C�/T��C<����!���:o��T�v�3R0`j�>��V阜��[���EU��J����dL/t��k,`��:RJ�B�I���'�9)�@j3VӘ��Jzxf���:��t�	��-(ȡ(�7�����#'�	�ÃɑBL��̞���z�CUr�ґ��˳�����Z��`��B�.�e��!������*�o�  ���P�p�.�
�G� ީ-F3_�\*TL#�� ��k��F����m��5����''v#S�5�O���I����U��1����m8�2g���j�,�dN̟����6A�2#&�/|Z:��VQ��7�y�$�I��Š�R%0�JV��m��x/�îع�5�US2*|:Lc��~8�e�q?������'*!�wi��b���B�rc��9�2�sd�n��u���KTH�N8�=��X��m�zݰ��L��5��=�C�7��8|%����>���#��a�s�_�|6O4���f�Eۡ�Lt(M6=��	�K�3 ˳��W �۵ω��
R���^8��TD�|Hˡ���r�����!i�,���h{�[��b���߬bOL����� ��]���E>Ϡ�8I<���Qa�V|�$!�R͆OZ�I���V���8�0�+&�ou��ӑ�*ƛ�X!�A����?�����ݹ�)�gY�d����Cn>�S�����h�?��(`��c��A�f�[j��2i^��ɴ-��Q�a�� :�"C�a�٩���>Ta#pA���Q�a�����v�[V���� ��NWK��a�:�*��Q��7��9gr���!����	T����.�����;W<zצ;��f�^�Ppb��f�G�?�݉��Qs̵ ��A,E�欽��>/vO H�b����Y����+�J���[�8"����$��v՚�|�R�纣m��v"�H�5����V��Uz�H��FR�.�!2.3�ol�f���6v�p�y�I'%����G�{ ��W�Q����O\�+���!�D��Q�cH��$�\��l�e`5��η��roJ���A3O��fX�9�ixά�k:t)@�K���r�v!����/RF�I��K��X��Z��E>	�����S���WvOAu��R�&rD�;:?F3�"�\+���9�ή-R����Bgq����1u�Oت����پ����$��G��	�5ۼv��I��s������E�/s����8>T�*L����]�#���{��̸��bM�~�N�5�{
:n��ll�\m-�5�����ő��}O_66Gxc��~�-�*F����, q�r��AbS��R�p�g �$(6�*B�P@fޢo��vf�_^�餻T�"��1P�L��9�O�tq�:��Ջ�������n�.��FA�]��q����%��-4Ǝ���	J-3���m[Ư;��0�k9���3e�ځ��P�� 5�cLю�S$J���f�N�!���s��_���
O�4���|:�ǰ� ����i��[o@"4d��8&���$�<�m�gh�{��)=���.�!�T�V����W���nz[sll��g@�g�Ȭutr*`���:�JɈ��g���7[��Y�?>�����1Ԍp�(Z^�~�^S8}�Na�HQɣ���X5k��Ǆ[�·��Z@�$�5�䲜�PGu}P\%-���J��c �j�
���Z�s�	#�8&���fWc=�cf�����#َ��[#��0e��	m&p�Jr�upL2x/qA������&T&��e��G���wQ
,�X-}D������Q��`k@��%�:+0c�
��s�$�M��,~��ɞtp�Ϗ�&�=��4p&��e�(?����(<��u���9��k�=۳'��hDADh�Y7Y���<yn���:�g�۳��]�i�`��#&L�h�<��<���tY���snm��rE՝KIڝqɦ[ۖ,�O=�e����W�}���\�\��XqU��4�����{���`�o�Y�3����sJ�~����KW�[,"�����y�<C�"���
ԅ*��+$f����h5���8�!���ؠ�D�m����o�+��{�(HwF�n��bFH���e�;������a��RRuS�vo�7PM�%��pF����0.��>W�<4s����I����@��C'�qæ�h~�:���a��Go��M�ݣ3�ߩ�-U��^�G� ㋦�~��݄FF��9jF��8U��F���,6q���O�ݙ�ƛ��l>�诲�Ȅ�)ka�M�Lc�˯P������K�!�r���S���k�6,���3��������F=}A�U�1���]��6Tʗ�U�0Q�ͧTԁ��[Ԣ�K��E���|b�~�٧��MTh�SG~t�2;0|q͒���I��X7�dP'�g�t�9��"�PW����M�;W��ո��QE�>�&
�z�Tϊ�h��*l��qi��HSL�r@�x��U�!����i�<�r��G˫ZBhPt7�Vf�4B#��`-�ց���
V�4G��c#X���,3|��k�+Z��:]|�GY{/�4<u����9W�����R�H�Oܙ����B�2��F'hG|Lԕ\Bv��q�e7�o����|�&z!�S�;�m�O�UMg�S,����ڮq���$��:��d���H����Y=1=7Y����Ls�6{Z�z���"���(��n�H��cӠ����@�j��PR�f�?g\dL�|],Y��fz�]�D}�����ch	�������
�)a�S���9o����n��%�|b��c#��}�t�&�q���e/��WI�oE�S��Y<��B��0j�zV]����y�mx���H�x��T�T>�)p'��$��N"�����=����2�Hp�$�v~�R���W��<�vP	~��	��ӭ����[�BL~=���f���R��ps�~�?���G\���P�V�vS���:j満��͚�'Z�ƖH	����UR��K� ���"��nd|���|��iӔQ|�2"TaF��|<�hZ�(Ҿ!�M#��n���v==Rky&P��G����}�
S�>TL���x�p�R^d3I��5U�rv��ڲ�K<o쑘�38ǼQi�1�������p�������iw=�� 7�x��:�	Ѓ�z� 4k[607����P�z����i�8���"��#F�ܓ�✐�����U�i޻"Q��f!6�#"ؠ�j�vհIgu��Z���@�ڟ ?&�}���;=���3���1Y�ɲ�n��v ��H����xN�g3��\>�kj ́�-�~'!�K���͉9a�Jp���_� d����:�萔�%�/D�]Tz�a��kGf�[�������ML\x���y-AN#b���R�OJ�8�9���)�4����d��"�����AO�.��@,�ni����&L�	Z�jݠc�ב�ϐ�G~j�
��xR�s.m��k����(����O�Q�ß`�"g���o:	�yF6���,A�����e����Z,\��W�����%�'�ׂS-�s�B���2�{��tƙ)���H�b-γ�E��&���`�����H-3�%�N,4�'��Ts�ȳRK�E$Z�q�[*4��
K����ɼ�Ƴ�* ��j��WG�WM�~B���6�mԍd&�9x��F�aO�"�]/���Ք��W2G�x�|�^i8h.CҪWl�c�����x{��F��dI��.����w�L�yr�f�'�M�xc�
u2�Z� j���5�qo��W]W��cIB�V��m��6���*4�r0�� ��f^��{�����A�l."ɉ	��V�?�Xj�