��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k����W�z�N��VXi^�p���d���e����}��O��_��؍ݝ�VI
��l�4��N���;���t�O�����,����C�anQ���GЄ�Y�<{l��,����%A�j����\e_�G�/:�N�՞S���}uf4���z7������ X[=��q&��W	]aA��?�g�c�����R���}%݆����J'N	�7�>�A��|��dUHh�GW���i�'�&fD�8�Hl ���"�1�D5	�qǛD~:̫Z@�6����⶗�_Θ��L���H�j;��W���'����\��}���#�<��-^=����Nc�	i��D�7Z}H��ʦ�)e�ϋ�{��V���Z9jL�X�]�JC�87DO�;��o$&��ޗ�(����Zvೋ�l7w 1Z�.Q��æ�����բ�|�����@����s�.!pH�W+CG���i���F%���������pk��&d�>�ɘ���,5�3����	�n�3�Z΁��T�
�~��q9�j��7.�8�U�I������Qɪ�.n���P �bS�).G�m�6_���2����hLY���j�	۹ 0������h�B�)�����䇶��t*Q3-�0��vt�L�!h�󏠇��%������w���b�x�69%��,�ݷ�������=�*��t��P��|i�M���I2����9O�N3s?��c� @�P��O�-}�2Z�-��2uf� 
"�Mz�gR�}���P*�X���oZI��W2^:E�];�F P��k8շ,<0V���1�"L+oKi�{�1&r3Q�]�x��]�;4���3LF���ͩ+��T�	Ϩ�=,�h�[׼Ғq��9����Kr(�M��jWe7�����Ɉ��w�4e5 .���e���͝��r@���C���zi|�rS�­���戮d��L���Hҿ�<_�<~����Y��7f�Ϗ�O�QMh�sj�:b��{G5�vA�:Յ�$��ù�4��,��ү>[��\��B��&J���ӟt6�6�O�UF	���{�^�MR��|9FNݽ�>�	:
��FJU�&Ω�]�|�^�-��i�޲/�jh�~�E��{���{p����7_������b?:�^	Eg-��g�٭7L~��?+H���=CI���_j�$[��e����5�eS��k*u�B�a�t+�n:�lP����0y����<5�R��?�=
�&�D��*�O�߼�`l���#��O��Z�pz�����yY,c �U�50XE�����q�S�_����{e2�����ϕ[�^��&��k�K�{@���F�&�����(�ս�ۼҰ�!��*{�]��2R6�[�3���ٶ~P[���pw�y#wob�Y#���0�iP����}o��q��Ŋr�h�-���\�l;�eY�k>��^mXgSN�3����ej� heQ����t����ÄuM�r@�.����G)cX��3�r������VEa�6�C�;��E����0���4ȷT����l��'vx({�k�$��^�.�O����pt�"���xL��õHL߇}��x�q��U3'�3MZ)Ww ��O�j��B,=5�	Uh�wۮx��$�*�L%�N�2���D\�eR�5;�\,� �^ܒG[(��=Wi�D�B��!.e�R�	�*���E`�5(YC8�d,����9�]p\���R��ƕ"��r�s�/�v/���;��a������U�m���?�jt�%S�^ �0�$��Qi|2"C}Sύg��H\߸�j��
h0 ����#v���@g�ɱ�)Y��!�:]%�@Zd!ugc��ݕLr��W���^ɐi�bm��3��;,)�*~z/��j(6|Pc �����ѾG�E~��#/5����Z$20�\,;@�9��}ȇ��;{��+լ�8%mFt<�]���t�f��QZ���oP?��S��<���:F�~cK��p���	6��1�����oi��-�m����刢�������8������ih�\Lê��~N��WB���7	G�8�d������q�ȡ�ۢ��ޒ}Y���?���d�Q��
�fc�ڨ�7��.M���ҧr� ��=��#�kV2���uM.��	oL���Ā�:�v�e�X�����) ���� ����NN��qd�|�H�>�y/F��0E�R7"a4Q�9pv�n&d��ذ�	�v-/@O�������tyт���3(9����D4x�Z��v��_y�ŋi�{m�u� �`��CH�nVy���c�"�q�,��B&�V��"�v��ߡ�MUS�kK�f��E``�9O���+BH�߯��^`���Ʀ��3Z
<p���2L��+���?l��)ր������v�H��dw����9rn��SZ@�B��+[���!�a�k�1J0����Lb��b��r����7,<A���ɡ;f?k�a��(Z��������7�qq����.��tp%��mL�/@x��5���ę4�Ť:��*��'5������t�%��Gmj��KN�x�A��S���<xC�}@
W�o�e[-���$9ê��D��������jR�@}��J�Ư�O�MrX�5v�'� i����t�n���2��K ��:~���%��r�� 5û�;��L�m�����M��#�]�]F�6j���������QH��1E��/���X�����ol"�����}��P�����&#�˫��p��u�gDq�U�:˿1;*E��@e����-/F���i�|W(�����'�)jN�[��Xh{e_0r�	�1;�y5�ws�n d�Y�;i+>�vw��^���n#���|iI�o�'\_U�>"O�U�D�{i��~��դ(�f�F�1�׳�<���{�@	ǲ'�Z�t�m4����!KԓN� /����<���	���6�k%��S^�3�ń ����+���x\;���L1&�C�����ƚh�E���Ϊ�]bs�r���Z�0�)�4xշU���Q�2j=�m b��ԽT���~r5��a%ݿ�L�{�����%"�߁��mhJ5?ڌ�������_xJ&������?Y�1s���9��dʐ��cs��
��t�	�����HF�ޛ�^��<�[�F�-m�rUp-z��4�o����3F����5����z𝋺p8{�9��<�7�.1Ϧ�Op�	���!-h�b!1i'��ӽ��H������9�ڡf�6��$%�!��:�.�X������X����6������^b���e�N�^}�e�"�>H��xr[���Y!ԅ�����@��5{h���AX~��F�MK]�[P�����B?&��lS��7тA���yfn\��a�s�:��7�E����)��:C��II�aE�tG,F����P�hm�|��=���}.��E��n5E�,��	�Vˀ��Va�����<�o�1��J��4�����5�!
ܛ+�r;2��������������_�&���~b�-�eyZ��º����Ѳ�f@�W{[Uh ��`	T|�����������=��Y-1���s�����a�ֹ�z���&1�9,