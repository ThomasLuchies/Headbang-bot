��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k����W�z�N��VXi^�p���d�����3X��#��¸�3%��O)���I�n�������:nA��+�js=����K���K?#�o?Bɼ��۬ai!�{*^'�%b�l}��($A<Jw�5�<�������/=��k�K�տ�B���K����ѝL���Ƙh�`+���&:&ې�t~u��N��M���R���*�9_!e�����σ)��D/���/,&&�����mB͝�U^��?��qK���%nF��x˦��<qu+w�'��Y��N�O�b����Èj�&����C�_�E�_�>ho	bC	�J��犒��8����U�Ȑڐ)yd¸H��41��5IUi��rz�Cw��{�Z�?2=C�Z�,��H͓���y�<��>�2���0ED����t��s�&YP?P�����g�6[A9�й�XB<��Dhs���Ĳ�d�W�.ơqa��mxk\� �����9B��W�ke��c5��1�иw��^1픽X�A	>v!����
��� q2a�R��[騍�ѳ�5�Pn�p��'%����S5rԇ���q�)�p�g6N����xV�.Z�*"���NZ�#�c	 C�� XǙ�m��颯�i|��ڬ�%��*���2�2���>�[l��@��$��g�9xw9�}q�=���)���^G"s�������󾳵��u��TpSP��u�d9w�kp���mX���!l�%7uJ�m�Gӯ��RLAH >���K�bNzayn��F}rQpR+���ϖ ��'�cA-������#b
�`���t��-�0�a�X^w����h���y��[�ɻ��w���o�>��؍V�-3%�,���pvA�����y`~���f��Nxa�y`~����p�I�z�`rNs��(G��4t�s�}�����tuZ��g���I�=����l',�E/���Y@$�Ѯ����&��]B���npQFt>6������������ߥ�[t���R	>毱f��ğ&����q��<1���ݘ a���h��HI�G�x2���)�\a���u��kx�?��XL&&�ٜ�j=��f,}�N<W��ȋ�E�S���j���qHv�K"<��(|�q�����>i�'ƠL�}+ϑ�Jc�0���Ԯ�{���࿨�ƻ���^=�j?��.�j��q��q�,e=,?��tץ��:��m�j\���,�sq�ԑ�&��C�/�R9�&(�Y=�>�5EbJ[�dP7Fc>���Mv�	Kv8�J��}�d�^;�E ��ɬ(Yj&��q��s&��K���?�ǖi�y��y��J��nYL�ZI��������0���7�lps�^�p�kɹ���rt�a���qf��=c�jw_�ё�et���٪@��'U�ț${����W�-���ER���e���~h��qv z�;ϡlj�D��u�!B�� �N�v�\R;�)RHW��t�¢�����Uؙ��ϛ��Ley���H�pٚs̚�U��T�舎�'�� Y�[dM
�uk�V�C�e�0f7Q@�MIHv�w���=�4&��7�v� B�+��.�7�M�[�e���`\[09v�
���P���ṕ�.$u��*&[5Xw9�fy�&v\KFa
�af��U�
�8�"8L�s4���9Cn�-�=�EI����7���E�W�CL�y1��{K�з��-a�<��}g}�:�PO�BS��Ԣ�W6�1�|u6;��Q�m����#K�������1�?o�T�>_=�0U�Uvw�Z,�)%��v�	��α�X[��i�hʤ��Y�t�`c��FD��30��da�Mv=�`4�4͍0����ΛM:쉠g��$j�{G�;|�6��0��� w�ݫDm��U�d�("sXq�����;�����!�n��̟�"�o/t���s��)xsp���O�:�����7��6EA����p�˰Ǐr\�&���F���Z2�u�B���SK	�;gt��)� �.����_�nߕW�=5f�`�����jM&?J�U���mb0u���A0�ӨJ�͎%U��z�E��/�r:G���^jT�ө�� �.8���(�������ȆX��f۞��k�a�N�G'v���������_����Xُ/��.qmƆ|	�(�][Jq�L���<��T�.X�zB�NK�ܤw����`�3OۦWO$u�Lv_ms�pto%���x�F������f]J%����\J��+��ÐRýJ�a�1'�,␼�9~�#w�]�">�|�h%�9Ɲ}j�IE��;w���b�=Ӑ��'uE���`ܿm5���/�j2��<m�k���W��#T�B����*��H63��J7����� /�Vh�$��P�:�z�M#	eu��j�~O�����0���Qy-4�:&^���m)6X.�o#tȩww�;�t�����=���*W59ܩ����1��=�0�i��Ĉ��o��c��_:�gG�ӓ<	â��}j��1/<�e\ip[������� �L����1~�1��W�G瓒�Ȧ�� s�
u��uۏ�t��L��n�(s��dS��6�{G��%j�pP���	�G��h�S e�l���'gUhb�����Gp�=��o��a*��t��	����V?t-���>�`����p�HQe���Wި�.Ɗ��K����Z.���r�؋dUJ�V]��]4c����*\s���!/�[��d�`��}8T<���1p�W��b�lH
����5p;m�ܝP"̠�nL|6���A;)Y5�;ul�̀�a�Ƴ�o���t�)�d����G��:s��'�G=�](���O��ؔ�D/:� ��R����=~�]�
>jV�[҄��2\F�� hW\TWW)��/Bm�CXD�����	Q�R��(���T�J@�z�R7�AE"�O����:\Y���,hŪ��r%�Z��������$�o����(R����yZP��Z��ӡ�ʝ��|�
�b�.�$��E����(f N�).ɧ��E��v�\s^�;@���#;��� Kcu)g�md�&�j�����R������ו+n��4��!�	���)��[t\I���%
\��+�|�z̑���x���ДMH_}��a�6��	+��Og��̭t���m�5�0u�s} Ϭ���T
E�^���Nf�W�+�/cz�����5�q�Ԃ�T�W��Xh��B� ���_�/J\�}����C!,�I�~9^P۝���=��c0Z�!ݏ��<��(�י�f�{0O�F�i|n�3(WĘ�I�=�'�wf�&�ob��s�6��|��y�޵��UM�W ��5���n��3�����A=����%_-l�_.P.�K�6k/'8���}��h��}��_$����3�K��77��L��7��ϒ��2'b�P3��`�6�% 
�UI�!��~)/�Ӈ9�.���Gm.Ml1�!!-f�}=�yCx5�"�(K\5�S��5�?%e�F��ְ1��>�Lq,Z�ղ������D�d_kӅ��fc
�%�"XA��!�ZJ�X��;xV>3O��s/���=� ��n�f�ap��%"�P�<A�| x����,k�A�f��4na,HpCG��g�
���CES��Yg	�W}&�㴠1B��*�� ?`���S7�(h�� *S�*�4;zf�Zӗ�j�3�C���i���:~~Z4$��s��ٲ�
���~���b-��(6�C�?����7�H�u5��f��˒&��^��UIE��>)V�#v�٭��޴
�"m�2�Nl�������ZA�b���^a�5��q%�u���!�KT|��!�w��n�ʂƽ�p��스�r��W��N5��4G��q�����md���ޡe��	�V������W%JA�}*�����]<U���y�$��hT����=ѹg���q�pV�\r�3W��'m��g��A݌o�x��O�I�K�lC�Rv�_֨Q˜�<*�h~�����O������$i�Rj&U[�5bv��q����q��I`b�����9�R���1j4:v�����/s�[
�a��.��E �W
��ܣH
d���1�����^�:�IXYi�bXE&���p���L���8g^���E��ޱfv'���?���m��ML̦Z\9VmE�3���緁բ���}p�6�~��� Q� ����d�*�CD�]�F�˴"n����D�,�E}4�R����w�{��J�!Mܧz��"w�2�X���%sP]���/$�L�ܜ �#�>,e`��4��aiDU�ͩ?	�����*����0�֦��
��Cvf�U�mƶQF�ir�#�o�Lu��o�3�x��Y��Gv�`1tя'�Fp!VP���\tG[u��zށ�7��f�,2^�u���aF����g���M5dS�q��}����q�0�w�)�۷��F�Q��W�!C�.��wj^���+��๦'�L���
�r�f�B.#�4pCK�i������ ��l�j�e1� �0j�~��ьh�W��V��)�Ԭ9�����<�w���אWD|�����ZD��h��ô�B_��6��S0�∅J���v1��}E�����u�^����2
��x�lH|a��pܱ���K'�>�y��wP�����<.���q*�j-	�S�o�gVy��H���pg`��S/���U5��E��'���-����U�c��$�3��D��x�BH� ��{� ��5l���aP���<�T�Gs�HZ��+b��!������~�S,w��%[=���p�����o�V�Ǡ�������ӎ���cg,W�"yDi8�������i���u��D�"=��
��O��H�syMw�y}ZМ@b?�k� 'usӉ<�^H<� ��Y�@S��?�R*�=���M\{���im�={�_���F3���DZ��:d��s=Yxo־��y��Ϫ� ��7��cq����}(Bȝ���5㔵(f���q����'���G �grH|��\g��>�ڊwg:�`��{����E�_|g�]?�Ў��{���wCօp�� �ȗ�
7�4ƕ��^�z����_�ȏ��!��YtE����j�3A��t�� o�rg�)o7�s����9�� ��W��Ӂ�:6er�2 3�V�����,��X+����Lei���m��<Y=R�Xմ�ǰ��J����EI��DcT�pl���(I��,���5��]�'K0
i*��A��H��?�VES�i���Ӧ�T�8J � ��/P?w?��57�qeS�X�M��GIVT[@S�i�8!��5����i��hR<9���
��e�r��>)��U�k�l�8#��2���.z�pMB�N��.:ř}�MBJX�B)�V8���N�(9!�ޣ���jܑM��8�Պ�"�s�lңO%AE�-�84C<X��vj�M���C�3IT6!(��uЧ\��W>���Nw(n�%@���U'�-�rэ��0�;�I+��#p���^�RqԻ����R'�R��*X�^�4Z>���ꪯ��'Z��@�.�T����	��*NZ��y�
*�[Z������IX!�ӭ����tA�\"�<��jc�k�J�I8t�7	a��h�?�eU�ӛ }A���jWT�}��
c�np��&*�_ a�ۊ�\��ʿ����Sd*@J7V%�&�	r�,����Y���M%!�>���.�`=��4��t��q�o�$Tc��g,�yYrwjÿ��u�� �ꗝe��Aê����;2�r�P:���b`t��A��:���J�p����oF;��R�tQ��_i��]c>�r
Ü�����}�U���pk���p-
Ӑٻ�֗%��@M���ٖ���w�x�8J��X��3�<ß����'8sJ��Y<��_�|��[q&��ۨwj�r��i���S5�����v�+�{��kU��NFx���TSj�2��L33� ��+D�W��_M5��B���'I���X�Xz�v��th׌��Sg[��,[<H�s<0d���Q��0h1T�R0,�z��{��YV_��s��Wi]%l.��V���ʀn��A}��f+\0���0�?h\��A�Fu�Lz�Պ&��Ԉ��f�� �}X��K����x���BӮd}!Iu�#xd���������o^�c#Ϡ��6YA�o?Q�F��#:27�v�1�,�QD�۞�����Z@��)��9�9OĳK�����y��Ss��X#%�g�rIeV�-���mUN���!���A���V�m�A�B����nU�L�q��N8��~��aj�c:���+9�1|�`��;�ț�#ظ3z�H��w�j�vK�>NT���;N���g����U�?�P�Ixy�z�ym�<cZ�� ��a]�#��uJ}?��Z^k�^��U��-�	�&r�����*�Z;���7�d��j3� ��<�!�p����1�%��'P�#�^�g6�[_b]n���>�}����oˮM~5��7�ҋ*���[iH�B$����Fk�����������'�߈.���{�	�J#h�����%yf���F!דh�|�\BW(t��u¢��-֐�S�~���G�k�� �L � Tn=̤^υT�iJ�����`o���`��P}��b��g�D˰�+FYɃ�S��_h�P�&�j(	�ˇ�F�a>�:h��3��K}��i� �w�TC�eyM����-[ 8x��B�fO4
���J ��j�J&��eǸ���:\�Bol��j�����~;�|z~������YL�X���Zb%�����yM��������_�V�:1b"�F���I@����T�iad'%�I;�{��}Ĕ�K��Ԓ#��
5���I���=
���*�s�QN��x^�Jo�O��9#��.�O!y�S'����l�]�sj������o�Kj%x{3�z����%J����"aΏ�ABA�����yb�
��l��Ad���kq������\�D5�M`�Dz���M�l& �
�y�	)|��d�� l͕��֬Q$��3u�`U!�".��b��s�7�;m�ts������* 	C��a��K��(�\� �����lb�܅9TD�5��"��5*gjqg�� !Sny���8����Fށ��m��M�C)����Z�V������H��wC�X�t�b�X&�1b{�^���?{�V~b@�S�	��Z$���'�!�fN�3'�ԞiO�y���8�|�0�=�A�Zo��q�HU�9��8i����A{2���-θ'9�e��/Z��"B���z<�w�S	*La;D�f~���?�ڐ����Š�lts�/���;����Ǆ�頶zCtG��ؽE�K���+YT�$
��(�GKq�
Kۜy�E��+�in�2|�TTMZUC�;t^���8_�0����5Œ�[	9�wcgxe2εw�������OA�Z�.�N��0|�%�d���U�
�K�h�TCs�q~�.��u��'�mpF���@�@��R����sH\ND�%e�3���9�ڟ���O_�����~�n�
�8XT�&\%��'��K RU"hL� x�ȵ"���)�J?�eo7o~B!�-�`ePM����&���4�஺9-_Y���b���"$�K6����ָ�M���T�w[|-zҺR0<��()E���r�:-b���N�K�_�~'�U�:��W����jB�&�E/l����=
0 L����,쐷p�����3ވH���6�#$��l�ߦ��S?a.(=h��c�>wQ&O�,�h�ؠ	�GH�ə+H���nQΞi��[&]'Rf�t'42bP��ea^��F�"�V(;E8��_�r�}��v9���1ƛta5�b]v_��|ע����M[�gmO�X��x�H���%�"�Z&�c-gl�S��d|q8r��a�Nu~4����aq���M9ry�ڞnjE�5@ug).xT��:ǎ�NN	1��N/$ Tm+�k��~�q�n�,�zrxQt�c���U�hc7^X����3��lm���زo����Z�a��ў�H�5k_�mP.a[G`xg+�^0O��$�q��ħt�	�p�����m��26!lx�p�8�b�v��VH����`d�_9t�{�G%X
�|�sH��`4��"��¹|��9��^,.�ڻ�7����`��tQf9�P�,�϶p�V��6�����?�-K1�D:�$#M�d�p���<Ұ�sC�p�~�,��v�w��\S��G�?f�a��"1%�	 ��hԟ��9H'������j��J��b� t�,{���"���m�K {Z��{U�d�F[��`S�8��ɠlU�be��1)��7R��q,��D��-�<k4O��N� +L����'�3��&����U����t�Aºx�<�����;�����H��o`�+gud'%]�<"\u�r��I>!L,����Ҙ+��J�{B5b�@ˮJ��b"�K<H�+� �J���V*��pS0[I��i��]�T����U�Ľ~�7����=�&&>�~]��DL�O��@��]��8A�e��錾���'`0�:��FW�㜹���w��v�c�N�О�+�aᷝ�{鐃���v&�r+9Ʃ��5��M!�.�Pa(��J������3>J׿�S��O�OvZ����ֻ��[�l�/C��4��*���=�s�J��>
�F%f��s6��H����<cg.�،�AdنѮG�|�cCV���եs����K���A�CTP�DIg��Xg���(�*�h������a4+�қ���7�b���:�iӄ���ϳ�+^�J��|%~�$:�v�2�~>p���g�#d���(�����9��2�H>ȴl�2�C���_(;����Ān�����G����H~��H��2�H(FƝ��&�Wm^����D9���
J���I�k�܏lsҥڏ���:�&�	�j�3���F��Ư�j�ډ���>F0�/�&�[�r�-��X��F.s`��aF�R�}(�1;�1e1��L�2��;����kV7f+�Paֽ����N�u2Kɓ���Tz�����r�-h�A1�KC����~l[Oւ �L��u�O�D=\�rF��7���.�ʏ ��X��C�� ��1!�r���檏9���*|Η:a�8�vtO��y{]�)�f*�tE%}�b?wͺV;����"��hMnh����@ϳ��Zʅ���[���9L�$�c����N��uAdM���M$�F,v&h��ůtm���>X��|���L�t��sk�
�It�\~��k��PD�\�&G�[�Ƚ��T�?f��)_�����(�J6-7㰗�U�o�3*V��)a���X�M�e�5�:���<(�128��bq=?�����XV  ��<A*��KZ��~Mb��b[���d���ϰ�ݜ�Z�>��#2y�Y'_��6����7���e��sƦ���<��(<ǆ�����,ݑ����毿G��u�}Ia�\�X�����1I4D�xժ�b���YV�ur��r;��pE�KC�v��m ��uZ,�u�=G�%)hB��s���0�>Z��2�����4R�i�l8 !�pxtp���K`OI��;�]=~�b�X�����~emW�r��r%	������2�8*	�. �!|`VVsB��
��b��U�}��䱠����;UB��XfVX�SU@���Q2�R��i����W����7�k��6�����s�5��w���sGC�ڸ跎;o��ڇ.���)N�44�Dɉ�Jt��l+?��W�DݳW��yo��;�\����r�K��D�O�F(�pWA# n�ݯ�����s���u�����2�G����d����3Zz)%���~N@b+=\���G��T? ��)z,�X��y�2�@Q�?�L�h�qq�΋�N��ܭ��иV
�~�������⚶��"3�ֲ�d���0�
�R�ʄ�8�~J���^�f���
/u����W��1t/	l8�0��ZP-�ȹ��h���9\��4߹��p
1tY�/vh56a�T��3��Z�K��v�O����$̗����-='۶�XHH�b�^/�(�8�Ǎ����rr�|o���بU�yH�T���
 �#X�Y
�a�q���Nx��"�#�Xd�A��X�X�zK�-�z�\�����Dn����,P���@Vmd������F����S�$��%,���V������'`����i12S+�r!{H��d�3�1>��g�	AK�g���5Z�i���L�'	�5�$�CZ��t����M��F�(CA�_����.~�#-hk��%:�E�����d<"�.o0�4�R�$R=<H��뙉(�	U�����7iKЧPVt��������h?����'h���K�H�N�Um释��Bx���#�&�a�86M��<��]R��OG����޻��k%k�1ȿ��2X�D��ܓ#���5�����j���u5R�@#�j�;V���κ����'"S ��0�&���ݩ	���G�:e��vI5�d�,��?j(PH���ir�T����}^�pN7<����O�9Y$k�x4�!]WP���1��⤥�?hf��Y��l7����5&6O��>�.&��������ҩ7�zc
�)�����  �S$��{uq	B�t�����>P)K��o��qG��zy�ߏޯ�O���)U��4q�8��-���Uu��#�kb3`�R Q|�6Q�"_ࡘS�?�i~�nl{�Je3�R����i{p�|��{@ag�V�_`(P�W�l�ʴQٻ�1��Mh���ݼj)5��eĵ6��Xn'�D7��)Z�*��;� ko��IE eqB�"��y(2'@���Y�}�4��VJ!���ڹ#���q���i���(E�
�A�턍���e(<�[�w�$R|� B��˻�����u�;d�d�G��l�g�&5�@�N���F9�3�*��מ��zt�H4W���3�{i;îX��RW�gR����]L)1̀�;��t�ɌS=�*��oW?�7Ɏ�G?1��T�:��f�ܬ*M��HSF5Tl��u��4�5v����:�����N���X�`��vGbX?���ڽ��! k
���ͥ�9SHVu��^��3�6�]c�j�ẋT�@���Ks��zL������_��5�%���Y�L��@9��| ty�������0u#�r4"��-X%��f6l���H�$?�쒕b1�8����4�wPk��M����'��.nI��Et��I�bqG$�����'������E����;e�z�G�)_:��!�H���c(S����S����fak�҃�N�R~t;��Α;om���������|�ԙ(����	�;�� ����g��I���HB�4�1W�P7���T��:s��hy�[�ɲ*��I�N���x�[��&�'�Y���͉Cu���󶹬��J���"��[t��֠�evBF�!D������"t�]��Nn��-��׹�����C��zGK��0IF�����6���7�%�������3JL��C~�<`��<�D�#?w�2@��P�V{/ؤk1]�`d���~N�h
�mͼ�8�����;���ޣV���%cyw�T�shu��po�^�v���cm��q �H�6ώ�W�[(�Z��/�C#��G���U$�Hw�c���5���:$��n�z�0�g�Y`J�6�+��oA��=��<��D:~�b��=-C�/��?�]j���^
#�_o��M�L��>�*����eD��)/8d��b�Ԍ���ƺ��>�MN���"e�������2�](�!VH��݅���dE3��Ѧ]����*O�#a�U	ί�N��7�}�2��l>l�9�z5�8Z�i�'���mA���R^L������2
�A��|	����a`4L�*Y���K/L��!�v����C�̷M�8�;�6õ2�qڠ�sǆC���&h!"�@3�������4,���+���/�Z cηz��j���ǡ�����E
T!h�g�!��`ә��eH9�V X�9��o{&S�1���&|[��b�ʤ�����J~5���K����h
�Y���؊���9��z��8&_�Uw_:Q2�\RxH�����c;5z����ܰ`�R�@���LoKcw�2V\)�V![���:�]]��S�\�U����p`�8!@��`D7�.��}*i�K� M7�1�\�+q�ˏ�E�I%� %�D�QU��_1�3�V�c�r���3�z'i!�:ݪj̍��s��?d�zu�LX �������A�@�T���K~�U�q'g{Vc5q�Ȃ�vD��q�3�.v�=�.�m�6=�����ڧ�.�w�|N��	�ҏ/,�r������!���z��|۬ YD@V%X�N+A��Wri�
������5���/�v3�#���7W�%p��'��ڡ��1|�/{������J���#�[��8lG�n|�@�-kۧ?
:]e�0�f_<��#e9�D�O;X�������yš�4U�D���U������mM�ѾkBO�
Z*�t��,�9���4�}�Y%�o���iֽ.1N�O� ju $������ė t�$�������<',��*�t���Z�����,M��2ڇ��Y�`��e?͆�<�je*bP�����CgVU�i���XmP��Z��ԩ)��m��>�({��S2�7�$��%/lʊ��B>�w�4�~Z�����G��c���_�-�]	E~7]��qN�VZ��䨽F� jv|��e)�oG#��$iG�:�̅J������9�J�F��k�f6�SR�%J�g�7����!ba�4#ʠ.�;�#�i�����K���^�,�9��ÿ�[�Й=83��ҽ̢�taV-�,��=���"z؛�t�i���T=c��V3�<��7���v6K��hZqC�Y@��rNm�I�U���Y �nެ��!l���,
���5���I����w��	%N�<6��˃��Ov(q�^���y5Hh�f�tyJ���I��9}�B����(��v�Z��/�����b.�܋������0�����);�Z�kT	ל���ӭ]	�mv��Q�5�;%tW�h�ݽO�m�Z̗�r
`�QR�a�rQ�ý����tb�>@l�gS�6(��M�5E�+�8h�^nQz�i���(�	y���]U�;��b��	�`�_AUY9�����B=-٠$d�K3{�@,?�	��0�� 죕ʇ�G.���ش+�br���C�8�˭�hˣc�geu��5o�Jn�H��5����.g:N1�b��j�Uq8J��v�5ݿD��U�]]!�#ݗs�g���t���������U\���\�9��"v���6]k<�Ү������ǅ&�P� y	�3������{6ٍa]�R�o���>�̪��L�	_��b8\��c�!���ͣdR�Hō9A�I}Q� �������	˰*u�_4���oZ�B����n�܈���M�:�zh*���{>��P0�?V{�Ⱦ%��m����>��[��k�Vv�4�1w�Y�p1�C�M:ȩ�H`��7��r&W�	0	�)�a��n�m�"���?�:F~��t:��Kn���c��7�h�z��O�7��������[ ��y�ݦyY�j���<��z	�w���a��X���)X��9ى �V�*خ�x����9��'�`�Z���v�Qـ�X�?��t�Q�Nh��l]v-��^��m�9ݡ���BG-@=Wa
;؃F`�cy��&�.jL%X�԰Dj�sG���{������������+��$��\	Ł�����
ft�R���
xu�6�=��-*��˶2��
o-X;�S��@�,�i�u��-�^ɶ�N��ɾE��˾Q �����Ѵ�\~�=m�����^~!���Tz�O	YFƆ�^�t�є�`�03;5}���Y�J�c"��:�G��Y��V��m)���b	�W����D(?ח�]��	�_G&����Ya�6��Y��/�}W�2Cy00S1�b�Om���x ��;}���Am�hE ¼�4��S�#���2�����o��͊x'ez@c�p���f'F�:$��Л��V�X���a2�<�������a��^�g?�nJ'������*y�k�h�EQ{�������ό��3u��as��.4H�鋻>��i1����y��<����Mf`W-��}xC��J�\m�L�0o1Eͼ�'���yx�㗓!1��6�e�\А߾猐+��۔�h[�V���9`jj���.����e�RU}X�K��n���5����vuð�S�ԫ�f�a�P��i����x����[�@����N䟺�o�3�yJ�e��󵊋�,�̓ʹI浽>g�*uz�ƺ��W@�����D��%fx�bD�|�N|8�$�sr��)�xQ�İ����)���C+STJ
x�m���1wnG0��-#���n
�'b��-�bB�wL%h��7i�1kcp0y������K\�)�[ʅ��>,9�	Gݤ �)�S���&�mԟ���2~�R��0����d[g�R���a��xgW��oY�����
=�b��g,%f����p�B��ݕ��5�O���VI�Ր$���9��s��a���(�nbw�׏_1���'
Yb�|1$�D��Zarno͐d���OIӍ9��L]�̢�c�YoJIysu�j���h�`�I�G��)9��'H�)ϒ6H_���O���y-�ba��y/hi�"c(3Q�_��f߸������B��L��;�;���:X�!R���;P|�@O�ۻ?����<y��u�7.υ���vz�����t��*�>�攉t|����-��7�"�U�ަ�,E7�d�)�=]�@��w�>O(%�~����[a�Z��ƶ$beD�k^���KR����!�:Pօ����=$�	�l�e��%=��(�4(���Ož[X;_G|cҰȥ��7������8���<�% ٝ� �l	���
IO1����2"ظ�0��H�R���m��\��'���Ծ`�<SUyot�`8u�o
>?W�8?S�L�J�'�	T�v��՘���=�ED����U��~����î:��mhz"z��V^�Pqڶִ!i�eGLʜ��^
Ts�:9�J�Q�G��&�
��d��%���CI�o:y;e�cF��#�3$ʙЗ��(�|��� ���[�	��"H�ºHM/�)����
罙h��e3�ܮ���s��g<3�s%Cat�Q��+�I[8u�i���z4㖏��*	*�� o@���'lϑ�Vo���cwm�A�i�;���a�#��U+,�j~Г_E*���s�h�ԟ[�[�fS�2�K�}���UH6��4` ����%s�5@���>u�F4�3.���T�+t[�f`:1�,:��aN�fF��}^Jک�Ҡ��Z���ʕ�Y�^��$cǐm��\#E�!�*�=�,4��Gଙb�3�F�dܼ D��-�x\ԇI`�5i��}4f5�'���,%H
�ڐ�N�wc��}�ҚT�L���!��́���$�ǟ�ͥf�sJ�9�o�~0�����;Gnw��u�h����(�.��� 	#M�����p�R�����O~��!Gr�_\|�$�;����J��T�����%�ԸO	=0,^����9'���w佀����]��S�G�z��4��AI����`�B�/+��x+fGܶ"��wh0�}�����L^Ջ��P �oQ>bb�n��m0c3mF�:FJ<
��YquE�ɰx�c�X?Z�k���s: �#\f쑞�4 �	5j��T��ͫ_�Z�z�j���$֦��bLj�(�;詍v����+:�HTU��2뷔dy�|���|Di�� A���}�Y��ȅX?T�ʊt���崚o���܅�t�Z�r�4S�*�'�k��`и޸|_]2�[w{�=p�q���Q9d�k�:8m�*G�Z�������^��n�w�g��"�f}�����<'��( Q 4�+��\Zm��� �t@s�k��bl�'���@��Z�q��&��h�������JAg�/��g}o�ޕ/��d|rX� e�m�qzpta,S=9:����Y���^���5��w9�p; ����~9���fm.7v4_6pWU6�1IHV����K�D��b<~N���R7�*�V��-j�Ѭ�*S��QZ����wvq�!�J�Lxզ���]| ��KkK����O��o�L.���,��xTړ�~Y�؉�����Ax����DoC��!�Qd��z�cH�ЪW0 �|XO���qrv�jR�Q���W�@7QNU���1}��,��ρ��^g�f�f�gQ��W������14��븹\�Rވ!�5�؊p��*�ż�[�Vn2ܜ�N�~ѭ��E2Q1�����C���+�r'�m��Y���0�a��lP�|e5=��6���(\�����D�W����:3Q���bۮ��X+��N��G���?@6��y�?	�R�in�r9C��w�j��v�8�F��Q�F*݊�|xqV�KP����eSx�I�w�Q���l�_Dɸ�F���J����p3q}��U]Z17��3�����۩u�
]R�_o-������8ЧR�ĥ�WZ�|�;Yw�ϛ�E��K/
�]��N��Ո���(A����!u/� m~ŞAu��lC�݅Q�F9��if\�h�1{��se���[dp"�X��^9";�m�qQv����[�~��FÊP����t-�������7r��=^�@t����Y��3�.���
��ctn���f��\���D�3l]̮���Gl�/0MLa���t�Iگ4�n{�W�U�4�ݶ�Ȋq�?"������J٭-�6��`�YoGf�K-$�k1�.8��:��u���4���tfd��JϾ:��Q9u�m�	���]�T�	o8���A�n�W�սHN�
YH>5 �**� &C�?�\��c�_b}X/
��Q{�9�g����b7}����O��`�3P�݉���KJ�	̧�����yR�5.o2��pG��j VAa����B�H�Da
m%Qey����|�f�����)%�a���kQ�����2����,DK�M����q����>~�i(o3��F1����G��֠%Uˑ�A@��8_V����8Q&�(s��=�*����]�O��ΊH�8���k� ��Ĕ�e�ykH�8$mM���?\�=8G�����vo#o�ީsلmG`
&��E9�~��?�EO<79�`��ӏ�iG������r�H��񹒸��}�k�ݣ�~�ww�_�lE[�udf��d�W���b_W6v��Jz�H��&F�=Sҵ!�P�&�;<
�̐����ms⻁��s{�J��_>@�ٳ
�X��$�=y��׀��"U12H�>~�y��{�,x�g�D62�=,�rq\���>S֢_�IK��B��>�Yr�)���F��[�a���_�ٴ���Q�|�^��ñS,�����防��sh���G~H}�[K�@ �i�{��q����"�Ov����P�_,]�s����g�j{�ky��8y�
�����g���(_��H��g���f�8$xow��F��aIW�&c�8�*����}ԧ扂��3ſ7}�oOg�c��+h-�m2U69����A����	�80T���!m���@ ��#2����A#�,���}��4�RU�b�<Ei/�;`�`��F����P��T�Y�R�֐�sH7٭7�� �SǻE^y}o��� oΡ7/��#9pԇۣ���D)��y	�t���xK:R����dڳ�"��s�hx4T��)z�,K��?�����l��n����@�s#>G\�*�V�ߨ�Zʊ��d1�f��Ei.=p�OSk��c��~Ú%z �	�d1�|�ֵ��r&����ZII�e�]Ŧ
���&(�޻ä˰�6��5XfiTF�Z~-nx�u�߿�F�=�V0�bo����)�r��t�$����/3�%c�z<��]�L�d�����3C��n�/4�:��d}�\~m!\��$j�d���ۄ�o�WЪ��_��$�"!fƞ!ЉԒB�9�M�/���6SH'���
����5Խ��н	+��K�؅�-M1�V�\xo��v��=V�8>`����;��9��r�P���p��lO�/e�ct.C`�O�+)��pDZ�|Q�L��@0X� +ti0��Z�#xUE�����[�I�x�o���M�t;��{����W���f���O7�Cݬ�̓�.эb��#�3,?S����\���d3�'?=l+`JAg��8`__�гpq��ࢇ���:G
��DL�������)��,���j>;m_�ܸo��^. z_]d�v�P�ⲭ��QM
��p�J�vkw�#'��R7�PU��M�,��O�+�����>���zM]�ϸ���,'p{�21�r����K�T<ͼ�r�:�I�������)��i{�c��'��N�L8˞���/2��\r2����;��G˃�<��d�Xں!��8�/�;B�b���0N4��Uf��A𗺃���u����3p���i{vv���Ǒ�7�ԄK��#�*1kX0��{1c�"��*~	�?�\ݸ2f�5a��8�Dۨ֨�U���T��>�k��(v]�� �-���3g���q7�����0�S�W�G`�bU���]����\��ɞ�[�w��ٽQ��I §y9g�˜ٿD�L���,-����U&�a��W�a��	���\vCz�?G8ŷ�a������KY���Hv��(�q��+a0��Q�U.�*t�%��^F��+��7��@f��]�Y�kq-N�L�C+���W7�qq�[8���2��Lz�7	�7�t�n��b���<m	��y�ӿ�j>�oyV��
X"h���@"�ՔId�ֈ~�����/}_��ɦ]��O['�⟂�#���e�#��>��z��7֧U�Yj*ҩ)��2�P�=3�`��-�KEC��T���&A��E/��7�m�ܚvn	�7��.��hla{��(�u�&�"�$��+é��8b�Y�����1-Xj�L� j���"���2�d��ʜ8�W*�Ql3�@o)����f.QH��������ǝϔI���YFϓά9G[SYO�������6�� ܭ��Ș��L��"3s ��(��APg߂h���E[ϱ�;"��:4,�ө�<�4�\��k1!��g��c`���`��B��Bݘy4�,}�#�Ю�i��s�;^c�wԝ,���Xx�]oFѿNb�t�/�-�2m�9։�ڞI�E�w,����G-N�Ӣ5�0�D��H��J�yH><z`��(���c�VwF�z�%�>�#/�-`y�(s��(�	%̰=}F~�:���)�Vx��`�\d��<G�iO\���V�4��do����o�0Ƀ�mj���?��me���	dn�pɏ[�,�	{1]}���m�%"Q��w������`I�ĘeѾ	�G���m0��A����i�Me5)ܰ󉟼�S� }�����J����ͻ�~ZRo��T�_L�/m�Y��΃c����:�!�V�8����s\J� \��؋�f��]�D�j���0�d�Ǣuz����vx����v�ÛL����`KO��e�E���A��E���T�} dl�1	 r$�k� őơ{��<o!h�{j*��Y�Mt����^*k+S��c{�d.�co[��j���n�u�`��rf��t��3(&/�˂�D�"�3�A����� +��A����W7@��^"�����%�M�]I�h�`�r�Nݘ�44ٓ�<�fQu;�a�J���>1����
��@#�P}�J�n�1��Ey�-<(�ך���ߦE�NNp���LTn�����`l䡧�e[�L�UBN%!��a>����)��:w�mv4S)D��2i&����{cO�9�hS���5@��^W��*���bGB�=m�Y�k/Zȿ��%M����=Xy�e����eY��d�<M�Ȗ�Pi��j��wvh�b�� ��ۊ�7S��e�LB�v&��,M�E��~��c�؜Cu��zp�t�~(��6ikOyua�qU&�����ED�x���idJ�C����}X_�ʓ*�K�2�2LY��J�(~S�����N[Hw�?��Qk�:a��u��F�� }��3ѕ͋,�(��7�C�t�ق.s6�^�4}i���fM�;V�����.�����,��1��p�X��N�`º��UrOJ�����I����G���	���_-!�y���l�޴�qN���W�(���L����"�ص�>�/��<`�Z11c�,���i7<�DC=�����2Hq�&��ĥ7��"�xP-�i����m5����?��xQK*;]f�FɒR�v�5�ՓʕO�K�lf_�Xw��<3��.��pE#�g"��o�>����v2s���*�u��7o�J��b���18���A����=z/t\�(��F8�Жu���?I ��[	~���᠓��9д��@+���zn�"��>�g��2hK�eV>���;�Pa��_�Zrd[K�uN��s�$?֏H���I|,�� t5�����R6s��'|QbC�F�T�P��Ű�M�m��؛����?�[��|�W��G�4 n]o:�~S{�����L��z���b�Dך]K&��qv���Z�5r�f/Y��� l^V ���ѹVJ4g�v��|�Ԏ+p��o�_e���T���t���}rw����c�)l<Q����ΩN���	�$�m,Q"0r�����/f����O?1Ǆg}&�[�%����ke��z� Kn����&��,��	�Ъ�
�gue;�8�����LX�CɅn�ُ���4�Œ�,�C��y�����]�1��/�������(^�����4^������P���a��ȭ�&p��%R�3�=a���r��E��#�Əs��p�a�  {
�hC.���0��
��hˉ���[Ln�<�Ӱz &���:#r��>JJ�14uŐ���OׂQ3-�������i��)�{��C�\(b�@&�܇3�Ă�����J!���u]�u����bǶ���;H(4۲�o׹S`��1�񊋊?�Q硷�������u 2���bR��<#���Z��$�����)�Ώ:B�dt��f��z�0Ӂ_���(�Nf��%7���тw��a����v!|�d_�.DZ�~�w��˥�������e��y��G���m_�n��oF��9�;lK������%VtzM��Ӯ��m�$���u#�sy7�*��'$�3MG�t��G�n�@k�U��w���ɳ��\�
� P�gzK�P�.Gדݚ>�=�M���SG�S����1l���J��$Zx�f�	U�>HRڌ��̲�P����GP4����a�Ѱm���7ǵʚ�?q�\���8� � ��%��幮dr$V�o"�8J�*,��ar��Ɏ��4R����V������zT��1��-H�~�v�c����߄�R��<eHNW�	��U���4,^'�>��$q�8D9"��]�j#q�C���`�������)�'�+�G�,�\�RS'�Y����M�b(X�?@��آ?�m��j�F�q������m�y���^�"��Er�/�E�1`�� mD����	��e����e�C���>)	H�(q�������MB"K�(��q[{w��ɕ׎|f�����1��궦Ë�q|v����%�/��?��(���)���Ej��w�0U��6����D�A �:l伉Q`/�"n��z5��T
#O�".��q���	�D�z�Ը�b����U	�؃D$�$)�!��K������b��Q[N��:Iy����[��1�n��^U�N������&M��)yb�'d;���oLJ�N�\�Q�T9��՝$�~��G?�a�	�FDtr�f�YXE��]�s��8d`}�t��,�����*�ɥ-0��`zv�������{xqi.a̒�-ԚM��p�|�Xs�0����D��k͛�ƀ<f�_Ct�6�fL�#2:@q�|N_�6{�}5A[~�е8�l�V*�톋��S�'�nG �z��@nOb��ri��I��׃dN/=d��/E�͠��'�A�<$�xJ
"D�l�Q���:���͎�*{���1lO�<+��-�p�����d*R'�e�i�cýQo�6E��Hlf\Uk�a��&�H�A�Bj.d� ר[�����1?��t *
����N|��]R[��ǫ'ɀY���v��=:��}��R����T,	��Z��k
�k3��y��T�}�!׸�p�M����݊t�F.�������㣫���N6&,�ڎ�T�E��C8<7���=_2���M&�Q��#y�4���+,�b�+Nf�u��j^}uebbZ`��(��I�2g�T�Y��V��g�ԏ9�����C;�D��B}.���Xx�F#g�V)4T̖8�EE1h1��a����9��p������U|�R�*�f��#��d�5W��^d��y�G�ϸ�t�zȳ ���*��w�U�H��7��<q�E�}$�ì�$��O�_c����MT��(� �E�d�q��pԓ�K�R%z�D����F�w�k�I���]&�k#��W� ��`>m�T^��h}�@�]%7\9#j�g�75���U;&,t,����[�#�MG�}��8:��J���}����<������tM|��!���D��d��blru�p�k)����U!ݔ��Oۿ�(�gQX �e�(t�L�H�S�Hv����$�_�^�G=�蝒u⯇eQ�J���2�=�����EWS�0� \Z�͋,��W*�j�.�W� ���I�n��ޣM+׎� �	�i-��ğ���	 P���(:��t� ���|d�*a��aD���[Y�X��L�˖};@� F��7�w��)�wB�q�ZuYF���`d0�A�r�Er�X��,	W0,��yfo Ȑ5�7��+!�iFr2h)��u4ƅS��H����� �i�,��+�%�6;�P���޲�7�.F�6����K�}
��"O�)�eك��^�<g�?D?��A�R݆N7v��1�@�7�@I��1*���Q��&פ���2������jH����xg��n7�MO=��׫ ��p�g�[?��OL1i��Ժ�;u����1䴲9�GiF�?�`d"�P�����K/x�eMa�o����)�@O��!arm� ��RZ����a�Ogd��v�O����+�a���s��\f���j��HIOq+�x^��Fʾk�\nE翂�n��?�>ϵS�s�� к���K��p��y�g�Ӡ�Mˉx��j�,0���{�'y8|7�8���'�F�[
�!k3s���4�Kvd0�H��д��1�RNU������G�'K�����<�j������R��k�WV���"��)^�x{������s��0�����*����=��`��
����8OV�����=���=PC�����^w���2��[pv� Ҡ��:�����ս��Nr=������&B��/�4�E�e�{���ۅ������"h^<8ꯒ.
�}�pFvv*�����ףe٬�IL��A=i �oz��w� 3^���8�p,A
v���=,��ݽܤ�����s���}kH㱛uw!;]�"��N��7c4�DQ��`fԉgCB�5r�m�3v��z;}P�&N;�����C��RP����6���h#1��ɮ��FU�0y��H���r�u���)�}H�M����]��:�Ϻڹ��x���Pn�Nq�0����ה�����WQQ)�0�-9
��y%ş��j�MS��݇�u<?q���q�;(�����Z]"
���'瘒~_����b���Lתw_���H�U��dYj�1�#>[��K��f� �����A�m��CM5��7�p�U�g�"1V��4펖o�J�,d��s̐�p���VQX�%���kƊ�4w�����G%��t@W~"~,n�&7z|2�|d�ʅhFY_/g`aMwb�e��`�F�&�� }�Rq�e� ��߾�R��.^�cS��;#���"�j�����0��F�$�4����^�����h���v�����cO�#T�u"�Eܦ�V|R�/�R����J3���gz4�T����\���R��x�W���Hݼ�����EIL>߻�އ�� ���������EGS���br�!2�.q� R�@�����TO����7� :���Ѣ>���� ��X!�L��7M�l�,���$q�
�{����_K�E�3"A��$悈��oԫ���>�ѷ�ř!�nŤ��a�e�Y�̈́En�ل&Q�{�p� ^	Cf+� �.� ��I�SEwý���7�`�[>n
��{IY,���Z0dL�����ߓ�V\��%#e�cܤ��{�	�W��(�7GJ������~�i$�Y��,�d7���Q�._�sK�SEn�D�r���!�3�
qխ��|��6��� ,���8�.�"8�`�_�9m]Հr�ݰ{T�0�P�9��?�--��z�>{L1�D��X=���_nл�H�|$�w�h��C���{�����d����+Q��L�Du.w�Q*f&xʐ�yQ`�ԧ�Šn1�>�{[�gZ*�-wU�m���|�X8]��ikOV	l%�J9�?>ف-d ��aǲ����:�܁���	��L��3����JiM��E����׈^6��RiAG�vv�ہ8%9�JΩ�`.!�f��mE�Anſ~���
!�(˖�1�`#k�!GL�����\F������6�j����A^"�Z	F�^�������D�Cl|�,/c~���C��nx/S����@�jfN�:y�� e�j���q
�Ԇe�a��c$�5V�zW�#���AՉ9_W�Ls o�h^oq���̙�~�_�=
��}[60��#�K�h,�H��YY+h��b	0��H�Qq����r
<� ����ue=l2lh�:�r*c=��m�HpY�kY�LP��=�@˽���]�hb9��4��WOo�,��II������K��u�ӌ�i�錣��!g�߅H�O�/y|QLh�>M�d�]g ��j)�I�V��E�NBDA�v�.0<��5 2v��Aư8�+����V���)N�SQ��(�,�������Z1Ā#��Yx*����C#DL�?G��l��D�v����)����;I�e<޲��
(���>rcӖ��A�3>z����L����n�N�I�n�鷻�(ؚ�����W��l������"A9̥W4��ݙ6a�z_�nd�{�)H�Y��"�ʩ�����`�a���<7��}����2�E3o ��5j��3Bݧ9m}�\�H�+W��I�!��pn��\����ebi�M���v#�NT�s(����m��b�1�%,,��`k\r
�l�z�{�U�P�� ��9͢�!���_D�-	c��O��{p3ē�r�W)�:�YTE��5g0�~$۶��s;��0f�sҬ����e��u���D���a�C�j���8��eLc��Űx���5�{����8.*H)7�փo�Ff�@2�MoE*e�:IH��	�?�bH�6��ro���'<a(6�y5�x�����V�1D�B��w�(x~p.�� ��e�zU��i�չ_����<�+�u�G3߰�v'n,���\��y,~Q�t|^^m龭�}U�7����Y�#�����s�G��đ��-�a�1Ϩ��&�f���H6���
"�`CY��IչT�����Zs$�
s1'� �V�2�j�`7B�Qar �t��{#�q�zuk����̽����U����L�7��vDڹ�ߥu��1�QH0ٴ�/c����O�."$&#o�9��F��3��œר����_ҖH�\Kq}�J|�Y���z�A��,�V�%阄����(� ����!�#L�f�s&����7n=���MY����&C4�Ұ�!5Ț�j�n�OJ���ڑ֩�gԉئ�~�\z�B�W�ox��De�I7>e��[!���z��S��("������eW΅c�/s/�v=��A��)]�ƙ�}�e�~t��xN̻]�Um�!�]����xc��ע_��~�pr��zz~��/��x�s:� �"JY}�'K@yMǇ������fO��U��B���PMĩ8Y����ʔ�2))�v%]d��Ρj0�ţȣ:!�;_$ >�󾪫���!�r�4��k��nCuW�dM�뫷���0���g_8Os��ͦ2�"�{[u?�Rm��j\��n�p�G�	X�gE�ҧ)�ӾA=��ʜϔIO�3�6��@���f�38�f�T���҆DGf@�