��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k����W�z�N��VXi^�p���d��� ([����UZ%Ø)\��U���'|�}��G �{�A���&�+�Z�%Tޱ��@�۟�E��@��9J
�5����b�G�wM;�y��x�_�男��m`h�gK��u���]3I!M`�T	-;_������Ѕ_[1x�5]�:\��χ�O��j�����;�kE�a��X��/0Ȟ����U��9(��8d˪M_��\��D��x3�F��,r,p=pE��ErA����+zj�� ����ġ���Ʃb.��/N�b��q��]�d�f��ʘ�,��Ѯk@'+��O4siΒf���e#$Z�}��Ǣ���-�x���L�2�N���+ X�(VZ�r��Fl�K���vҶ��a\�=�-�w�#���~O���֬QfE���fS��K��q�#�Dh����.��V�'��`�&`�Z6yR�}]�RS�˂����G���\���s���ǂ�B+�AƂW3�/ēH�:��'eFE!�*��sт���)�=��(����4�
�cgF�"���{+�ğA� �/�#���I�V$cvv�����g"<�u��(/Τ|O�oON㫗X��g��َvm��;�Gw�?r�f>��<� ��&7;���=M��K�X�>C���j�&#�,>�\��@��wO.��4�40����sA�>�n��i�b �Ro��VTs*�M".;�F�_��;���E��,��<��q��}:�H���
7_�]����K<嚋��t �_ħ��2�<Tr��q+}�/Gi�1�H�4-yELC�m�3(CX���[�/#nT�2��Q�j�+E���r�y�F�{�x������y�y7��ho�,f�HsU����J��DE�V���7R�b�5��sJɻ�8���yI�R�2�KFiC)��í���R�A�������!�f��k3��]g��� َ�|.7EY7�e��M�򁷖V,�H�5�Q*S��'�
�e���`�X�}���Qy�����a�fOw�3cU)�KCs"|��B��s�����:1ڭra�=W���I���M��?5��ϼu^�SС!x����<��.k�u �]JS�T�j�nz]��B��4n��;��^��|~�_bM��]T�?�!F6����	�tX����,�������V_B�}�CCB[@�L!;0�a{�xZ���Q�L��_�y�/K�[��V���)U{���o� ]�K�����٨����\k[�lP#Z�������oJ�oߚ��xa�I��܃f����=c�R�Yӫa�ϥ:�us�u��N9���{їf��tw���Z��4������5W�OuM��[�
���V���H&�Ủ��q�0s�����F+͵cP�2�I��g��b�g*�}�K]~E����/�Ej͍�I 3T����&8f���ԒБs_�(���@&�M3��4rH�%�Z���'U�F�y�V�5&�J��ˢ,Tq8jx0F�r�C�0]��*��D\nO��@78���Dh�I�����*~���pt�4P�4l�'��).����Q�d�<�]��C��ೕ�c&�W�i���z�bM��I��y<��~��H�0;����dI���W��S4{��!��<0�Tu���k\�k�i�RCG�Fm�,qT�3�1KYM-R Fk��$��d����8
�>�j�m��]X��I~. ����.��F�0*O&�;�I�zo��B���%��C.Ⓠ%�7��]X��˕A>w��8�>q�T{ �M��}��	�"�ҰDdO��n�C=j�vC���3�W��+����:Q;�t]��C�]��2l:��iN�1�܃�l"��� ��ku�lo��z����$��4�g��H��[�{.�.�����ۙ���������`�J|=PS�a���(�[�R���+�9��$����i�p��	4|/��� ��!��h����!�V9&%E	���q.�oS�x�)[�5� :#�}�o����ϳ��u
o�lGZ��ϭ��F#4�H�H�J�'��BZ�L��*\[Bq�'����|�8LRo���a�g�����Oç���p�vJ��i�x=3ֳ(�i]Z�v�;����ղ3�+Ҿ��_�]H:}�#�ۯi���bv͒�#�O��4�SMz9��; ���,��.̤�-X�� �fܕ�+~5��I�l��?�Hi���۾鐣�󽮢w�2qZ`�L%M>���1UE���Q���E4�9ѥ�!3�GV�SHk
y��m1X�f�Q��2w1���8o�
@t"�<��D�� !=teգm����oJ���̊��z/�q�����B�5����sȫ�.Z����$�Q�(���#괩`����1L���W�k���3P໻��r� _սmhs���̹��,o^�*S�m��k�,��K<I�pO��~���I��(+��Lc�e�M;����V c; ��{k���x1�z�dMS�V�R���G����?�����fR8�hbU��j�r��ϱ�/v�ӵ�b���¾U����\�b��r��l��-:���V�6��duX�8�QI��%�q��� ����Uग�4h��Z�|
�9���WR� [a'ZǼ��B��FI�n#�D>�
Q��u�ԭb��bJ���q�o�Y*��1�	;v��*A��ۃ^1�H��;��B�ǫ��#P=�^���f&n�|��3\�b�; �Q`�|��һ$�(�\%��O���E$��!�.{TMu\�&l����z���cU9�9ZY��锾�6�rj�D��9c��M�#8 q0��*����bM�E�(=�=((!R�O��m���aZCE$�\g�#�ý��]S�4�T5V;i��X�%���G�	+�G���8�{�Ҟ
z5}���"/�+`�����V���3^��ہ����-55�c^�N�=�MBv6{�S�7Ŀ��[-�VA����p�)�_�piv��H�T=���wU���z��o�xN,���d;�	ќ�_���W�gX}��pQ��Bp^pQ_[hG��W��EO�y��@��V��S���'��1��������o{���W� �>s�	l&$��բ=N������k.�g�b#��j#w$v��K��j��"ڒ�H���<��c656k��[���&_��!HGl�n�SG�~7ˡ�.7dG�ό"��Ls����&1�/b����n1����7GZ����!����(� �F=$8.��G^\
�Ri�HѬ:K:PYBE�����~����XD1U<�����]�Q�4�ɴ1�b��aye�
~G���@3n.�:O���`�Dw�s��g���4_��Zc�	ؓ�5NwW���%ea��V�I�z����\~�gA��H�SA9�uO7
�P�[�� ���ߨ�?M�d�|05�
p����2�&���3�y%17i���T�(±+�m�'��#7E7��@Z|��N�� ��[#S��� ���pm� �W�{�ކ��EV�Q�L��̻��g���9�\Ⅸʕ�LI�����y�Q��L�a$��P0`.�\�|��y��(��)���J8��������yD��O	�R���n
2���˔	T�J�����^t��"(K������<(����'����LcD/AXgN96�Ϯ_��D������i@���4�)�.9�aI�M��	�)��!p"k�unI��-vN�.�wmo�����7��n���*�ψ��b�P��>�`2�$�����/YR��6`�| 
�^�t�{�a�!���/�&��P5�C1q����aꆃ�14^�5�ACs	X{��܏�*�D���K����)u��~��ͅ���Yq� �\����-qa!i4���B����9�u7�M�Q3��ip���(�Q�P�Ӯ(����)w~M��]�^o6�}!\V��
~P�&)h����@���e�#p�X���7�Ox�%1�EQ�ф�J�6X��l�9q��ߐ\^u�cS�`�%̶�"��F��	ћb�=��'B�������h�-��]�D�F� ��͉�i1���Z�d��y'���Mpt��N=@ݥ��L����	tp$�%r~&-JW����V��Ǎ̮�=��G�^�#u����N����k�V<^��Y(V�ᡫ�'6=��@W��pɅp�;���U�d��\Z*�����((Y�e�z��L��S%�=�(�X�(0�OMn�{�/�`��
��YH*<�m������5��҂У��VnrZ	��S������䠷�&�}������#�f6q�[��%"L�؍����@�G�53��a�c�ɮ���|���n�h���G�2�}��T>=�����.�Tx����J���~� ����pq�s5
v����A�m�tHu��i��5l�-�h��y43U��~���*�Q�3M["�	]���~���^��d��%�17��ׇ_���5Ҿ�s��g�a�So;��|8~@�[0R�۲規��u�{�T��O��j���}�	�
pZ`f���
�r���~�33s)�Mg2���F�x�0H%%`�X��۱q��p�#��	�Ң�Wju(��_]z|�>�]��[W��_�Lx�8��2��~�Fb=��ߝ|�\!x߁�Z����<����cU���㪱�w�z�K)�����p�i��^�rWm!�5���m�%��?��"��|+��i������,��꟞����DQ��C��g�,�7r/=S(;y�ʔwh;W��C�SҞ�8O�i��{���G�'���mDR5�����cg�ãi���j�^D���Pp��?Xq���ÈT�Πv�)/��R� �t��h��`�e�3(ѻ�����n�F�Z�Ǔ3�F`U��?�^��"�2��]�ov�mY���8����Gq�;�b�!��0�ZDg��MT VeKn�}�S)��!W"[��9�]�z�6��jC���V1	� �?|���5:�j�����^j�ì�j;-��?��aӕ������-l����J���������#b��ɕ��c���LlZ����R(��S�AXyt��r�G�X�J5x0��t�x�<���	�į�m7Ņ��O�H�f��_F9Z��9�g&�,�i�6R��(���?��t����,���v���1u�:	1D��< �.	rk��G�&f�Q��E�,+Y�����)�S���g�s{�md��Ȫ}$r��)Mt�	P���qq��<Д�3H�>��A+u	m����ˇ?���3p��yXP[�