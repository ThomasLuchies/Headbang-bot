��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k����W�z�N��VXi^�p���d�����ҋ����C2F�
�Z��>"�.�y,<;;�I�Oۙkء���x{�B�O3��0Q�Dy����I�p��1#C���޼�}��>��RvŴXH="QK��!����r4�K�"��o2��	��� ��*�xP���]�)RP$��?N�a*��Ȍ��[����B�:��T�B�}��ѭ���K����lM<%l��%��U��՗/7��ȗ�' m��-X��Xߡ*�զ�t�wm	�⿃&�4bgў�w}Jh�&ˋs���{���rX\~d x���ҭ9ލc����/wA;�lq Q���K��Z#�SWK�Ȏ��PHח�撕�Cj�_��Jwp�H	��np����]�.��f�ع���rK�Ͱ�,�g|x�V�b&Le�F+lMv�\KoЂf$
�~�Fj��#?[C��0���1L��mƗAB4�Sf�@���� �,4LB���Y*sT�Z���q��P�Z�j6,���r�@��0AX0�>�l��s/�����khx�nZ� �e'���fydĮnĪ\b��O��6K࢐=�/ �[e�����_�"sG*]�k2�����f�w�]��5Ř�r�g���٫�z�U�ZL�'h8#�̣٘����e�Bxb]Q`�Ǭ@\+��d��
$n�.��(ف���$Ź�����X�J?/�Uc����:�|����ri�צ���������*��	��V�t��5��{��HG�:����&nx���������������h8Ͼ�;��\k�fA�� ��T�1?�7�� �m����79Q��s�B�z}g2�B�����}4�C���,+�;Y����R�Y�U��ԃJ�8��%[p������T����UX9�[Q��{�{�M�m�Y��/x+t��4������u��s��[��k��w1��C͂�e@B�d�~�&H2�P7@]��O�G�~:���G�S���g���͕>	�yk���͍���U�d�4��Uf��r�,����F�{3Q|�B$#(W���D'��N+3�W�+mU'UE�̢O��������b���(8)A��z�&�������`.����'���Sᵴ5���&�q{�J�M�"@�'�}�hS>BQx�uNY���;�n���0o2��6��.���gJ�!���r����� �{��b.�j9y�ӠXj2p(V
�%v�a�|zs�뒅%K�ۗ�~6`-���@-ȓ�
8(�;�����vH�����R���"8Vx��C��W��8U��e��d��bY�O'4�9򰠁ʛo�z���M��l_e8�w�S��uK^��n�&�"�))�H}��-�Y�'���8��}�0, �g�.���������8�PЩ98	<�ԥ��K�:P>b�@խ�����R�,��DE���U���Ӥ��xd,��VXR+H��,�U�v�G�y�^F`5x͟=�|���l6���IM�vc,��e���w��.�-�n����K99�V�}��q�ɀ�n&(x�c{��m�����Jh}hB��:�d�n�dIʡ�w�����{$�8Q 5��.�/�`�|z��Y�n~f��oAym�T:����즢6!3�;|�N¬
��ES�*���р�vL��d46��J��c҂ �hj~�P
���Dm��g��HWRU(0/�������N����bb�e �L)����V���b�˖��;��3�Z�j�ϲ6���As�q�z���몳�q�d��[���u%F/��s���TBx"�&�[X��Ep~�𜪫�>�p�!��YhHG���j?����<�"��י���-8𘝀ִR��u��39�r������RhQ�\�]ez.5���1�N� �P^%,���U4��  �||�����O�+��Xt���~�ھ�6'��E��8��H�����X�p�� ׳�ap-W�b{��\���kJ"G��7��/��������������F�d�t�KW����-�Jb��Km]�|P�*�Z^dL�Q���,Ax�p~��	�I"bO�l��3�m)����8��ѿ�S����5O���ג����a���8���g������KiǠ��Dc26���ap����0����&u��F�gO��k�Q��z��~vE�	1�_��r4>����+и�O9��� U (�B�u��/���c������4� y����8T` ��@��ڥNpZle���ޫ����-�@ �������[���{����ԉ��k+�c�5|=���|_Ln&�$ *M࡛�e�����8��u14Ue��\��rC�Z08�4�����k�Ċj��s!-acPH�>R@��;N8,��/�k2n<c��ҡ�"���a�x�(� 1E`���~a#���A��(���E�
��"�p$L�g�v��c�mY�&�sW�++0����b�@$�,�6Y�ʞ"���ů���gv�y߀��2�D��gzߖx���v^�8��|]_8�HZd9�ir�'%Q�.ߌ���<��H�jh�P.�h�w����7�%�.�~`�	���_:�#4�)����U6�{q�QO8����*�J��u+@��I7���]j΄�XJ��Z�uV���"
f2�Þk��Yd�(�yԱ�ؗ�'=F�踯!��
.JZK��(�)@�N=Z�rhhǗ�:��&�/>V�MK�yt�0T�����~��[�V�y|�<;�n�g@�Z �I�B?�Cotb8�1��c���	��f
%.��0��p俤�)�1k�V/B������>�X����"��ap,�R�ްA���.��4饧%g`G*,\9��J�a�hR%^Y���6WǊ�w��m��<#����7���g����J�p3{��P��')ǜ��?�K6�k�o)�(�ԁ�{�r
"��fѝːc�Vy=1�QlY/��=;��ζ$y�&���d&��$���ר��Z��f�?�ӿڭ�.z�J���
z��X:�,"����zV�wC�>�0����U��~�� �����({��T<����i[��*�C<�(ɬQ�#[f��7>�@LX�Q#P
��0�4l�X���?oO�I�Q�C�IUm�Ƚq] ��2��S���QQu>�n.y)�.PQ1�P�ngJt�C�SC/⻣>�$�
�Kf�"���s�����Y�69�˝��+;��W�H�9?�\ %�l=�(mp$}
C��/�F�q���ϊwj �CF��wq�y��3��:�T`E���6#��K���J��C�u��O���<A�M�.�wA�hz�k����2��5�+���)�^"��1�cw]��<����� �6K\,�ձdtR 	Ӟ�R�*)5��V�y�æ #	F��g�Wv�鵠�w�������C�5Nʡ���"i�G-��b�+��(�F:�f�c��+)�9���j��1e�'c�m| I)U��d}�%��H���v��v83��+�h����)��Y�·9�hڭ��`������S/�Ơ����P^�{��(�eR��/1�0Z*VI>L��d��M*ʎ�ԍ���0)�ڔw;���˂�x���Ved���+���P�T[�IkjЫ�� 2��i o�hѺ^vrhs[~�IۨZ�3?6A�����f_��?p���-Ճ�͑R:1%��(�x<��F�"��|TP�ޞC���給Ie���%�8s���i�;�[����&�|w	0�@��q+��� �Wb�9.&�=�X訡��0��3�oI'!�ȱN��2�q"�rkٓ�ܜ�-[ p:$�����9���:-|�b?��v]�>ˎ��DG4)�9��) ���Ç�϶	X����,A�Q��w�Rآ����]�n�� �Z�_o�:���^�]�{�i\���:�W�è\��y�_�+��%�k_���JoMmn>�ퟛ/5�D,3�g&�m�NC�+ւ���K���'3��+v5���oH���'��t+>��m9�����b�Z�%��s�A�h�!�A��q�A������\$p�K@1�mח������r�T�.�ш���=��g��d&g:B>3�rh���m ����<֖�z�ʆ��a�Z�Uk��Y]��=K�(M�D���H��nGn(���sN�V+]�'�F^r��يK�m�]-5��ͅ���K�����qs%�C��r�CO9T���V[�)K�E{Z��\�,"YrY��3�z�?���8/j�V
6�e�%�!��~K���)~����T?@����(��y7�����5�������n�#!|�~�}䯿�O��
�1�����P��ȕV��/ávn����^�.>U4���ޕE�KDh;�<��7ÄuH����6�|�גu�t�y�)�?><8��ϗ=��>�7 ŭX���z��u�Il1S(���r�5%�Gc���F�i���lګ�b�S{B�}l"\�x�π��XU�A��s �������u�L9޴h�MB��\~�)B�1S&��&.wĭ P�f�IuZ��H�1ZP\� ΀�
:��õXi;	��%Ή��r	컝a���-���!�M��{U��aj.���z���˱G;��$g����#J#��A��zb�=�������O/ ����z�p�"x�ғ#�ӻ�zC��P��=i8�l~!����%�U��Heۭ rw�o�lK��b\6�PC���P �57.c��&V)pf��eN����~�4
:��7/W�Eи%5��+��fKB^����+0�t��h��&��;�3�B��@�s��܏%vF�P������d�D�.��w�f�����m#�&����6�]c*�c!?��Yש��F�����N�ְ��|�>�i]�j51BQW�\"\��G�4�mC��m�(%8�/O�x;ܻ8j�#��j����� ��}���r�|�V�R=f���o�@T2r���7��O�  �c�/hY���Zf��3ν��#eӥ�_��$B@�Ng7�=@������$�<�ܩ�.�I�;?N�r���E˙4u�#���Qi��'ˋ-���BP��x$����I�p��P�:C�X�\��k?��WG��{�;�IC�)'�ZƦ^r;.��әj�0�����y�G=5�4��F�d��Gj´���%ͼ�$pi��eHe�fh2a��gÙ%�J�R�� �I�5a�����v�+g��kJ8��
�V,��Q&�K��ˇ����ʮ�3_�b&(Z&�ղ���p��/X���!Q_u՛�n��MT�kK�r2�v�F��	����EU�CV.M��Z�Fw��7?(O;]':P�V;��1��e��Ѡ��^:�M�������v�,M�8�qpծ�<���w��Y۶M�6���*у�����Z���WU�g������:�R�ÜfE��]���7�1Y�=�k7zM��V$�҇����#�[���n���������:�:e���@����#)q,H�,�n�&�qH��hF�b3��t�Òm���f����q;�N�L�bø2���&������;�x��"f�Zc�M��k1�9q�$_�(�ː4�X|@�=h)��x8	��X�a,D(b�M�|EN��
S?��b�ᚸ�HO��p~�2yw���S� �NI_z~��,u��e^.0�&���D��>ɭ����?�+&��Fm�&T�]Kz��$�!�Ņg�����v�k5�T���\WȚ��+e�HŅ���g8��/�g��u��&�ǫ��]�]�E��h� c0�����3E�צ�H5���9��ª1�����C��^ޙ�=�c�x�O֓�B,I�>x�"�.U+���K��{�����,;އ�H�
R��_ǐ��	�>(a(Ə\��L��I@�Z�+�i�������>�����̑|�,�����<4!����=I�1�b���޽��`�}�q	�����-�+�'4�Ǟ��Ƴ~aA���7���a;j�J��7j�!y�MK9����%o�tk{��Q��^�>A[������ΟL�f��U<d�v���Š�Z�s��]�(���NR3�Ѐ����2{�z;ǁR�f藃�-�Ӻ7�����kP.cNn�&u	�+)�%� 1���[��NQ�|�*�TDK�k����ܫ����qR:r��q��.
�{�4t�q��
>DSl�vP�)Q:y����9܆L�O���zAv�`�I1*r|���N�o����^�I�eߺ��9F��!�~��Y`&���~-P�{=.���;>|	�b��+�����*6b�u;�u���T�����b�N+�'$��kk�pV�`9q'���XӺ��]������ڻ���,M�ֈ�b�8��ư��Fv]����6�S�mw�?!�������V�'�5B�_E:]�g��aeW��[���Y���۔�-#A���������ֺI���U���e��G���gjO9��	��S��R^�xS��f�Լ`��A>r����d��f<(�٘�h��w߬y�=�zkd�S�������x���$�41����Y��.�m������2�Ɗ�����72h"�mh#�4+>�P[�k�,�R��u-D�]�R��v��1a�{j�y\���D6�A'��,�h�e����f"$&-q��5��lR
;�Q�gJL;�iT�F�������C��[��9�yF���Br�z� �?<�\��(Y��f�����H�Ԛ�)��>eE�r�p����#ߜ��j �.Qc�hL��Tdm^.M ��v��,���s����	z�?!s|U����(7ujo�0#�������-\VCm1r��w��UpN��-���"�[�Jƾ�̞G��,�- ~f��FK�v�#�(Y(�v�L|��*P�vj���ޑӅ�<��`[δKk|�6c���-�\!p���x:�i���
��/?�y�=�q���
e�;s��-x��AՂ�Зegd I�C.=�[����Ha��	��%��d��)W4f�ѭ�#��-�s\b�E�ю�X$�K�4�qh�\K�F{�22s�z;oN�y��t�巏|������y.�_txx�5%� h�{O������q�j{}��5g���T�l�L�����~[����o��B��J5Ҟ�Ik��5E����d� nBŞ�'~�E�?a�Tb�Ѻ���J4p��c�u��@?�?��*���e���G{�#$80u�[�a(����n����ե�苸I�)ƴ��?�`�}E���	?F	�?���_���-���J���:� �Mz�gH��2?qu�0�g	>Y�����)IJ�IV{T6d_=�A0�\�+�QN�wݪlQ�/��Y{,���?B��8�����Qp�u�ɔ`�*�Q���d}3d�YU8�wM�Ό��^���P������	�z�^��������p�3���"�������6�~yy;�W싆��QK
���#���C��S�e��v5�d{��%/��6�\�M-�����{�ն��2����ƻY�QO���χ̢p��m_:	�A����͎���D֥RQt��ǃV��UU%�Ǵ�!�Tϗ�;��m�[�<oTg
��|����cP��k��=��D^��)z� ��v�y�1-����k���S]��"���LE \�"�1�Dd��%�+��w5!�=g�?�h�6�����@� ��$R�
��,po�)>K�n�8�]���:L`�&��}�#D�Z)Ŵ��Xe��r��,��#������}��fw�D���(��.��w4B"p�o�6��'w�K�w��rW�qW(8F�csr��!����.�+���=�Jn�J�vOw�)�C7ž?q�@��������]���y��X$pG�����R�	���)ʲ����[��A����dٰ4��g�N��z,Fp�����q���6�Ub$�u�&���&�֒�3���>H[7�&���ybJBQ	σ8շJ_�ʶ�l5`2L�/��N��ӏN�B�v�3Ҙ]��� �`L�v����U�䓨M��5��fCb��sw:&z�=��K��r;|�m*-�Vd�t)�uQ�GqUo���w�l��ؐE/h,�ؾ��i��a�*1cM��i��;S?
D�z�e��2ѝ�w �X:Gv�2�_�ۑ�i��d����~������{m�IK���7v:g͂č���u.���=�rذ7�5�/�s��C��la������������ƞ�*��������x=�1�zh|�3C�[$`@�,A��b&Y"�R&���%i��W��A"9����s7�K[�̸@	}?P��lb���k���O�y�0������$�&4�I��J>��X���nP��a4�L9oy�(�5���I/q�N�[��Zb�7���m���A`
X�/u��&6J�zɍʴh�7����U=%p�,�����Ce��?�j�5�_"���y*ݴ�2�����q�?���;q�5W���>
v�V�l����KKz��#k�q����L��H����2�9�i��~9ޘ��~�e�������M�d�@�*܇�	),-?h4�CF=���w!����1���A�/�%�{�ω��ݾ���[�q���������:1$�t��ۅ�h�0N�}K�e*Ԩ��ؼ�-��[i=+ĲY�:BR��㮷%���$�(W�s�R��o���͐V��[��i"J��.�
���\YBC<��	����y���/�o���{����.ڒ�����&���
���H�UĮ�.R���Ɯ������n)�V��'�嬬�d�#�Ƈd�5w�>���������f�XzRS���)
�c���s���C�~t��5���	Bч$0��3�K���~���:�}(K�Z�Q)�H���!�w�I�L]�7�3�#`�Ҫ�J=�m� ���_L�ãK9����4�QnQ�w���ա��/@����ruR�,?An�Cl�<��Qq4�sol0�L�	k6AͶ�R׫4���S�n�~��o ��D�����>���f����F�M���[4�0E��7��Xh�VӠQ8s�����8 �I��˺�9�[>�W1	f�st,�guuoOM���7���AW���W[fc�gԿd[�)S�u�n���^���a��0:~�K��K��U�G����NuHYqc?�;ĭ�fQ!��kr�&7LvR��%a���IQ/���űϬ�X�>��銠I ��8;�M9��y��>P�B,-=Z_/��zm���̓����<B��ף�|ċi1�6�����vL& ��1�m�n����$�gF�nOo���������6O������񟴅J�[)I��Q�#��|T�j����3���]M��CI1I���u����ؑEwیs�C��N��	��e˞K�d������~���^��T�P0qO�w�q&�*�����z��B�ެfO?��9`�����I�t�.�HO����{=� H5�d��� ю{��̶���-�/����m�3m����#�!0����7��o	��om��U��Q�f'mM<M�Ʒ0��)K�ߗ���7f�����l��O�I_�éU/?o�Ob'�v��;OH�
s��6���j�,DJ��o�:�E	������,9.+k[T#n�����Kq�B���!���^0e�*4�֕lHG�B *�|����X�����j�:�p�!F��;*N�MS{Z�������y��O���P�,���<�<�s��o�P�b~�prj�Иu���oi�	��0����u������,�FkB�4b�s[s�������_C��^����<�)P�����Q�:�|^!�C��a' ;_��f�X:S\~U<�9,J�-�����z�c��n{)d�|@��[�����Ml,�.%$S�>
��)�G4�Z>���.�'�ف�i����d0w]����Ll��ꋈ��T�0�g �>�:璤'�I�*A�=��6�� m(N![Ǜ��i�{)���c���� V��倯�0]���G�-�?f������2-A)�����|3���6 d�|�xf���Q���i����l���嚞�C�Ǆ�5�Hl���eL�;㞌�{��अ���� ����o=f���Zv�b���B+���2�Y� �J�E:[��L���?>������\d����{��:g*E���$q�_�Lq�$��k�Z�zJ:��+�@%\f#
�;�Y���*wQ`OyiM����jB�"��ZnG6���Tb����]ô���x��C	_�L��~-dc��o��B�X��]�Bb�ѽtĒy��R�+.$��{��V���i�]����n<p�������d����Zx�G� ,5a�Z�e�� C�1���#D��?��/��Y`�VK6J�&�Y'C�6����B���*�W�g0S-����p"�Q��T�q"<��k�{�m�Z��K�_}�U�n�ք%�'���i-3:Z:Ů��>kN�|��0	Bof˔�.:{�+�͑F��ONw�#�}������&�>V�`�4$�F�q��gG>���=p�3(+|{.��i���qRbH���\j>8��h�H�Z#�X�A�k�!�M*��b�u�E�\^����Sv	�|V���m��n���l=H��߀�N�C�Sfn?I�P	YaE����&��n��ZJ�B�O�fn�j �_��X�Z�?�m�.W��J���)t�)jxJI/�ͳ*�ܛN��]v�4��9#^��?`Z�gG�q��%ṕWh{�H��Ӂ��Z��M��� ��qݶ3�jo���`G��{p,8��|tޮ)�T�7Т���͂�[�bW�N�jl�������4�ͻ[\hA�S��Ot���ly��YD�o��}ٸ���1Pd�%���W�Sjr�"5�&�A��2�XH���[���$%�LQ^�ϯ��B�%��Ћ';�����q�W�w��q�BO�ڸ]��<����F=U�0�Gp�!F���M(�P��-HhS��S@�v�U"^6fsQ:D���k���������$c2���Ǖ�w)�]��%�Ƙ	��;�&(+�u��J�z�Ԇ�
ߣ�׮�U�_���K���e�U�~��r$�UI����`�Ņ�G��/�ޣ��
w��_�3��j��$�̐��q�4�̯��<-�z�U�o@$Z�x/��1�b�-�a�x�z�i���5)�x�B3���p�/�*7h�O+~3��3�)��G<^�k�j���ЕO:�T/A8���k�HZU��d!z�)aA֯�U	n"�7�}ʻ���QU����pD�_B���T
OZ��#i�e�WE��Cz��a���4;۞0夼ѓU�kk����Vq[�����M�\˰�4�c3�X�P��:�f׷f~ �)#��C��64��|�ЪS�o,�~Ft��»_f'��ķ��Mr��B�n` ,��T�����ý��P��{�E��V���/�2�M#A9$&�=X��w������ށ܆�������3S'�<�v���[��8��d�K%F���������[A���|�aW�\���9�t�ɏ���,0� ���  Q����Oyc��P�2к7�X��dEՐ��L^��E�Fj���1os�����ޜ�����"���?�v-��FZ���$��Wk_'Z�OGP����؟ͧ��[��@�����8�_�����>ukb�S؅�,�����9�e�&
RKjxoZ/�_8�pF�B�E.��rBI�ۄ��y��ދ@PMhpH��BO�~P�U:��m�t�rgZg��_9dW�۫�P�d����C�}v�� bo.��$�C�%����XU/������uO�x���`��z��4��m�Eq�t��#0@#//�8��i�~	��W�?���
|pZD��.&��81��n��M�2��`YYB&�@�}T;+�����t(\I�D��o�'[�"�5� �!u觃^`���"�����Ef��<�� � [���'�"�wcp�5}{ :NG.fzWM?�%m��۾�K�LlM�ΡL�&V-�0r}�	^LH�P[X:�i�p=�j>���;�m���^�(��!��[����xỤVp@�H9��{��@ ��<XC�g�A;K��٨��%�u�]ra&�,�������5�H��1�E-w)��;�.�[��M��.td��-��ç��zQ����ś
��k����mE�B*���du~� |�����V�@f\����U8>�[����d�7��R>E&��k�0��6�����>0����
�g�1H�@38�Z����ߎ�B?.�Y�����)�ڡ܄+���e�u��d*g	AyK+P=b^2iQG�Znt��ÆS�οdm{��A��߱țt�ހ�n����I��k��3
�	:��n}����KDS��ɿ������j"���J�|=8���-=��A�+i��ml���Z�NPE�FR�f�:��QB���E�m�'�RD��ɯ���-��{�f�e��ଠ���6�b�άV	��U�!zd�p�����2���۲~��7��������=��p$����R��d��*yvF�xS���4R����?S������o7�S�p&H	��J� ��I#��"T�͇���C�\Y��X��\��7��p
��)���i�A ��]��ϥ9��f���oq�� ��D8��q�d1B��A�Nr�@)�����ӟK����:B����Y��n��+�-�?ݮ:�N����	G�{nŶh|�C��H>y��_w?PGѧ�?���2.��=���[�n��
�C*D�@�.]�xca{�ȪDL���Օ?�]Zٞ��O���jP���\?Tl��v�����X�2>��u�S�%��T�j�мZ���)l�=�e����'6��Vi�n ���p��N�,#�8�tTZMh(Rd�ٔ�q¤�D�+b�p���
���ӵ�J3/��0\V=$j��sBA��D{�?{ ����|���\g��D�2T���h˼Z!���`�&+����F/2�x|�A �څ�T��s��(q��g�a��H7L��{��9#<6bIc+��^��Ǯ�C&@����xy����3�F?4��"<{�yC��l�H>�x��gP=�J��A\ �S_5G�Р�s&9�y��߭�]�[�GFF�T�����m(�,�bF�9�2D�>�PBB	���2;&��^�y:���B�h��r�]VRt1E�mi-���D+��0?ͤ�[$�ˇyC�[�fIa���t>��ﱟ5_?����C�2�,��[
��;�6dչY<��c��B��EV�D��� s|���j	mF��_���tb�17��G��o��SllS4 ���<�gW�).� n�DHeT��7�YlQ��'f�ժ�#�
8��B�u�@�K��M�oB�����N�]�C�����0�r�2�x�\��f�y&��ߟ?�uc8�k]���U������I��w3����z��3�H�k6Q�4����.�_����gy�alv�o_666�V�m�-bWG
�ֱ��9m.����]��eX����׌�
.%.����h�==�����ȡ?�ߔ�o�6F��f�=B����Gb ��ߺ�: �;����>�e��:uְa�΂_��Р����V�*l�����%�s;��e���[��<8�Ak�L�����A$�B�9�;]�#�)��U�w�5�u�1RR��G��������;Ճ�^Oٻ�wA)���v���%?�ޒ�Af�%�@ɧ�د�� ��ѥh� �r�$b�%��Q�2��� �N�Z]4Y����_��oz�����j,�1	�*����)J�nP[�!�	Vnr�u3��Nz~W��_�\ިY8�0u(��i/��2B>q �g�ZN�/3�2��ۛ��ñ�Tq�";Ps��Rk��tԓp~�rE��0	kv������G�JN����K����h���6.}��g��
����/�arP��o ]��	^5r�Є�4��6σ��|+։�/�O1&V��� N��8�L$#��x��J|W���F�_�F���ͭ��@A��1G��M�U�ˈ���mtɂ�&�8y�4l�-=83*��*<%x�k������y(��b�,�b���S~��<r�2�H�]��x�`z�9�5"ķp���k��� -Ԁ�U��o��6��s+�o�2�㦌���V#�
��l�Q��Q��
f'QSR��2L~�RK�L���S�ˑ���;vcTe���������v�AtBHvv6�\+�`�û	$"�%�
�3�-�>31��v#��\$��� @���D�٫�)}*qd} �D�sU�貖��u�:�4YİtML�^'!��=�N�^&%���7��Re�V٘uf ��7߮E��j�L�65=�x��r�hnatZʯ]�rƸ����/恕����V*�򊞚q��A���i�Gz�D�����۰�0�[+��U�򽍁{���[�,�!VA��*�Xbg��W �F̅%1��k>��B��>y��M�B#�k�DͲ./�S\��Տ�I6���Mo�0��x����j�i*M䭍��`��Vz�x�O�b�ᲃ!��F�5\�кt���P�a����{����'rg�1�v��v+�������FW�K�}����EBw�D	d���@�aaC�V�J�Wdk�D`���i��u~go$5wx���E���*�l������!:G51�cW:[����ץ.�^0d(��}4�7�4Sf��V^r���E��T�'�j�C���s8r���#��V`rG�crB���	%$vz�_i/�vؕ��+����zE�Q�b�@��p���3��:+t7�S�H�ԇ.����"!���W{��lK!5��|�')���{r��G���7�"�3�4.ړ��#���(�E��P�Ö������b�����n��N��=�F�±u�7=�$"�_����k���W�T�j�[����>���w/ꏚGZ���G~RwG����į1$�;zI.R���>��&�D�� ���B1S&1�K�Ge����`�Z��`��ra���ѝV��Ћ�L�x�SEO*n�i���`,�O�_��c'Dꥡ����� �A�{Nn�vs���k�>JP;i�܅��ڣ�=���w���F>�LH�1&�o�w�]p�N�fXaO��t�|���	_���äu����'��mY�����_�7@g򖧋��J�v�r���p��+~M��������Ʊ�h��`ܿ*�`����!Ҏ�G��r"=�����ɖ��Gq�u�;�����Ӏ�0⺌�u��iqu�>��r�%�c3����g˹���*��aO0w	�
��PC���$�L�o��w�-nMў�燻8<+,�i�����' �����A�`0��m�ο�6p.|��3��$	����م/�/	�_��E< ��s��i�W���?}��J�ߴ�������oyV�i�a�����ˉ��2^���Ɲ�̳�����:k�̀���w���e�B�6Uǋ���/�J;�|�l&9Z�R+�$�����؊�e��Ϻ�㈆��/�T\�q�G���W�֏7�M���6g<��TwC;�ȿ������|/�'��-ǧ7?������ɔ-���ݓ�ȼ��%�1F��l��7t�-�/�C|U%�VDXN�DL�#�K
w�V�J�������R#�RO����é�B���v@/4�`3����V��
���:W�����U�B����j���/�l�?���C�� F"����cZs�zx`Z\�J�=m��Ú�]��C�z�Nq�*Xp},���yrZ1{�ю�
-�]�%������T�ϲY~^���V�Bi���҅�-�B�5^��ֲ�����sO�D4c�J��쎲�{y��o	�3���i��sp����,p���=��a2���@h�J���B�T��ȺD)�麨��?�ӓ�:�%�U���^�`�.�����̶8:W��9�} ߿�i��A�涤�"6G��#4DvF{D�͑&������қ(��xL�J�r��/���7>�~�Z~�Z�QiV�G����.F�ɛ� ��9fy����j�B����A$�	I�[�N�7tT�m�#Y�ʌ�}s0�d�*��ӕƥ�T�� !�[���� (��4��ד���C�&���~0�Sׯ����Tӂ�2p�"� p A�@�"�a��.�é�as��u�Z(9���{`�S@���O�=��z�m~?�����W���� Uo��e"
J�B�ks�Ew���F�����#6{B%ş���G��DzcE�E�7�A�QjU3ʮ*��	f��5M�f�;��e>
�:>�)�+ 8�}��&@'v���#�9�$E��z�����!@��R7���Nw�d���ÛAgϊ
 �}[uP���+ ����C�y�v����H�4ў|{<Q��.8�e��~�,=�� �H�p�#�w^���o9N*�`���M���y�%�}D��� )�K�s��F+ڞ&e��=\�x������!f�~��*b����ޛL���+IgK��+-�h|�J%�@��#ޒ�,�j1��;>�4?C7�s�)R�(�>;'��v�조���Fe)�&G�m����K�Q��w�����8az8�Ţ�P�]v#W�ى�� B�)�d/���k� ����z�ey	7e�#���m{�y��5��m��M(���>�N�Vp����B����S��.�}�;�,���j�(���f��CM$,:
3�CʛL ������?U��O�M��;C6�[g�>w�+�����jElg��>�S̫,b��U~�_�dL�A��qIR6�\x6X��G�"Q���|뚢��QJe�(H���?�_#׽���u6��)II��~/�A��Phg;'[	���v��;��T�D���WoI+B��*=�e�F��P ��}��8��A(��)�lx.���NX��TI�V'� /��ޝ�9�?�M �bo��e��qU?�N���A��˼���=�b�.���4S�G��~����oS��+\'�/O��f��6.����<a>V��R�l9I����lkk��3�;�,��8�;f���	8��q�xyB��~��2�1�}3bˏ����I&��־h*0�5��05&���c ��\P��mēK�#���<I�0Μ#M$;�ٙ���T���5!�O��n&5���gN�²xj5��ʾ����ƥ2^�k1����NS������OI���y�+�x�at�w�~U�gQ[�FXE�=<��$�M��?Yv٠�N5���{v!�Č�^�	��_��tK���M�`�q��*�O�r�뫰ƅw�xC���F���N����7��"Z������ԸB��ެ���3)�E�yp�.�nV)oi��j���]9��!��eX¿g����v��K��֩�O>�;!َ����7h|�;t��F;��\e|bX��Q���o���i�0r��k�.T�X?4�io&�HH��k�rCf�~��o�T�7�_�:��vT��G�+���jQ2����l���������	����ݑ$7��)c�㽧'w���y�v�	��]��
�Hß~��z'�٠��5��`i]	�f����k]�gm��FJ�ɏF��n��\(z���\)BtVX
̫�C��![����rr��r�~ko��z��_�Z�>;��$�ulw�n��X���U�D���lv���Gg�ġg�G�\���-���@�6�&���	�dO��L�/:��άa�Ig<,�A���xD��"���0��������
���uά�I6?<ߜs2��+ ���9����pڗq/{�[�%�6�D���I�fX�V���vt0���>=t'	Ջ ������n�Aس�@;`$2���U�"�E}�K�p�����3+�������{�I��;7�T���k�~� ��cl $�s���i�!��������5x�i����eMЅ�c}�۫��ͥD>�\ő��2�F��]��ݍ�1Ԉ=!E���ɉmR�qmj�x�%*A�j^4�x�<�krV�w����f(�h
��� ������z=Ӝ���`�}����"-���7��T�z]�$��Ѻ*�ss�/ m����fgy˅tw��D	U"��%k���G���$�҈��x�eB���z	�t��-��*������� &�oTP���FCw�-`����_f}|�w���N��"�=���J��Gk�;'�<\B���nu����������a��Zr��a�ukT������#j����ˎ��E�p���[o���+Ib�=�|�6����F�S@�O��Ȧ|asͻㆰ�m�!�Ě��h�0�v���P4��݆̐��jDs���ug��? �V�u���K���l���:} '�z���<`�w$~���	�Vc���N�W�-�G�oy����w�����ְ��.vQ&c�N�Ry�7B���iD�j�|�
�F|�~`J#�������a6���@��3����~��y=����U�\%�6~� (��}^��K��Is��wY��ĝ5���qB�!��lT�����h �jqU�.1	Y��.�x�V/P��L�� M(hj�Wu��>�|�a�i�SC�}�z�?Fj��Rﲷ�(�$���5���k��9R���н�8օ4aĐ��=Ն0�����j(o�-t�� ��/}�:1��Ib
�W�'�$栢֐e%�����Ľ^xH����q�}��!��P��9^qy&0�'�jZ"du�f�T������K'�Fmu���󥑤c�f�I�ҷ�5���/R���Qf�L$y���5c8~���zo�ݶλR�2W!+��'�p�jO Z���$�n|�
a��F(�y����;�3��pxV��*�_P��g�5R ������pU�e��V����ڢ#��!��{�������}�����%:��%�"���r��T�b᫩ӷ��|t�gM�}/�x���u�!@5�MqQ�yO�9#��d �j�	�q�������u���YD�f����{�Z�7��d0�2A�K_@��w"����W'�)'���a��UC8C�C,�U�V�7h`'c��(k�l�5�B�{�D��·� ��(�
��� �cV����2��M��"�Ǥ�5��I`��1*�$���q�m�1�b	�S�^��9o�>�0�r�D$L��ۇ���M�#���ϒ_��(Z@�J��-�S|��*������{�K�(F�u�/�~��m���0.��3����?��k�1�c���&uW���*���;\�w7�������sk����у������颂!%(.%�<_/�c~J�׫
������J�dmq
��W��VjJ��|���{��P^f�͘���,̃&1)�@ñO�E�~����<���oS�;X�'EA�j*���ޢ���]6.�\�ȁ�dХ1� ��y�d�D� ���L$��dh�V�,���#���٬Te�T�\�VT���Hb����ۀ��sQ�����?D��P��r#|+$x��c|j`����}t�j���{�E�ӭx����	r��"�N��Aڕ��|*�B�V�5��Ji�T�&�w�8]�Z(�U�o�Ã��~C_������W��{�[��_6_�&�4��
�m�:=9��MνC�&3ۡAK�P�w����Bl��3)�e&�y�.��8�:��2oڈ��q�8ѮN�χ����H\�'�����ztR{c�b���XF��b�c ��'�C2`g"�B�5�t�IPF���|��ÕB��O?
�(�1v����2Aj�9�QD%�ܘ=���y�d񋨲\0�o���d�b֝7��,+���X�L��x����k�� ���/=xdW:�g&��':�!���ZKj����DO8E���P�y�}�(g��M,#�u�Z�eNJьu5.�S�9�U���	����j����L�<�^ʨ�t�]S�}:��@C�i�;Ȉ�tt|xĿ�����Kʹ�{�Ֆsg�;�D+mI�H�c�ڋvPH���nu�J�r�zY�C�C!q $� բ&�.9�r�;y� �]l��F@G/�����T�֋�Ec��{Eʛ�zH}��O��,a� �s3�@���L~Mܾ!�a�Ig�0��ZY����N]*�t���'4��C
4 �;�E���]�Cj\T=%�A+ID!0đ��~���K-�H�AvIDې���l���eV'�쒗��5#��ύ����DZon&�����h����3�g�P���:���j��Q"�3X�m���#I3x���h2�K�pilL#���¡癕ϽyT
�@���O�����'�%�hS���A ⁮�%g�^;���O�3%���l����8���X}Z����@巊��L�.�q��}Q�=�RF���`p�].�|�]��s�9!�%�!�f5 ��$=w�ʩb�Ap!ЦgA��:���t�K��<��%���b�Fi����ZD&h����:r��l���3�s�'��d&�k�=D�rg�;l��M�t�L��D�^s�l��Ƭ�0E�u;�����R�űi\o_��%z�P7O�̶��"@�v�x Ft�GXRͦ�w���.е��#1).�GRƊ�/�	�X���م����U��������0>��ƽ��3��@!0���B?F�:_��x�B|e<����4�	ˇ
I��I��V<ݏ�G�wn�����)9�dz]\o�d/�2��i	��-Vdi�^:ts�N�b�0��������B�fT����T/tD�d�7��;I�}f�~�����&���̖��������6�SM6^�?��pi9�"���#�T��^\;�u��u��� ����q�1p��W�餆t���|,��y�{}l��w�������\��N�Qn��䯦��|�������5�A;V�sd�G��r2�dF�ڲ����q1`($�/��q�/.�{'�BH�#)�3��vPi���~�� ���%�1%�����v�C��N\�|m��
���L^��e�^Y�X�M���^p	Q8Ƴ��[�6Q�<��
N�N-��nv��g[�ƘG4���պ��7�d�����XX����jE���7[�[�w�]͘�%�����ՖQ2M��t��]V��Z�������9�����q�փ����-W��*�z�9�X(�b�:)��8z��