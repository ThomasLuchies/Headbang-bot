��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+�������;���ȹ�v{2� ۝ߎ#�W�ӂ����ݠ��>_g5���t͉□K2���Ec�ſ��`\_��cW��Y���NB��*�!�#-/�����0�����e	�.ZDG����g/G�lз������s�VS�]��	�_,��ܳЅ2꩙Ō��M=룯+�&HfUk�@��%��.���cm���pZ�^�&]C��l�QQ���UicM���*�qz��ZU�^u]�2�=>���J��מ�#�^Ķ���l�\*l^���F��A��N�QI�������T�xĞ��pǚ z���4��)�7�z�wcl9du�f,u���� OK���ي�H�I� ��l��.O � F�		�,& �����ͽ�`� 7�(������,\��S�!�4��ݮW���l@����1`q�f�>�U�g��E�����a�md������N���+���+���}���t�
I��-�&���I;c�C&�Q�J���5땕�?�Z|D�YP��e�|*���#܉B,��S�(����L���͙�p�&d�d�d;B�Hᨷ�ǻ��qa�+���  YEɃ��)=��������Hr߈�/G�S�>������`0&	�wu^+�#C)H�C��f�k��U�lv��v��״KOgC�Ѯx��X���8�xh��]�
�J\:�68i���Z�O	G���[s�B:�E�6M�x=	��Y�hw�946�֊0�緪&�td����q��)6��xK��BkWG:I��h<m���'&�4�>wz��5�1�)�r{a���l�p�I��A��mӔl1����R�GJ���a�[&ĉ���<¹zum��;�{��3s�m�a]d�6�l�OiP��k;PZuU���zx�+E&��\I��s�MD���� (���P�ᇂ����'�����	�6�h2F왜����[Z�F��>)�������n�����|e�&����'F����=��A
�ETj6٩ 7.$��ZYC!9��V���w#�O��a�s�q�W�XM��r!��x��|<1�m~T�Dּ��$�JcG�rl��zZG1ܔ�'�= ��-����$���&�_v���Y
��!cvk�@s)�zp4[|��%$��$�n'�v`�7k�����F�S�:pHiY~��UzyX�έB��y��D*C�D_2�ꆌng^��n��D�yI�*L���L�D_�f�Jq��EJ�ӝ3�t���E�]���<+͢�_De;����j &�i�涯���

zk8MX Q�?��P��M��?�4��`Z���F)S`�0J+��؃�K�=�����X�*�q��zVpt� q@`�!�`��1έ@�{k7<u^1+�[�o&�S�ճ�LJa��L�3A�]8��[n�)�`4�>�S�%G���Il�Ӧ�{���6jm����Y�H��d\$�W:D ��q��Q`�s�/­�g,{�Ó��5��R]}Ls��>�=��j0������q_o��ps�9'5K+��;Q>�x� ��\�9�&��E
Q�_'IL�T�a��	�#�-f��E�gG�iV���,YZ��
�bkZdF����'�@��i�X�OM�<��sjQ���#$s�a%K�_��P|��Wֻ�Kj��x���'�`3?�G^h���H��e\ί��A����#|Ki�%S�?�TB��7�GiH���f�l7m�-L���/��J���Zd\k:����ک�?��F�ȳ"�`8�ЕZ��7"Ǆ�+��a5��Q�� ���z���!@1T�=Ju��\��'V�^i�OB���*��>��;�T�G!�2f� �e��
��}d���F���6n&��|��/�V�GM��2�ě��;�]B�Bi�Ϥ�2ޟ��%	e$6C�y\ȡ��9"�kί��m�CL���Gj�X/�� ���F�3�~�$$k�~���'��齻�����O��<�)
��.� �$��k�ɫ�@9���yu��Z�c�ODk����:�v�?����<F|��d����|m��d�V�N��Ǎ�C[��A"�8tȐ��=�$��'���2X�����,��[�9`�=�?W� ᲆ�u��k��{{�E�yv]��\���`�3����r���=�1r���F�������n`����Q3~R���Y��}Bl fHN��G�Lh����7x��� ���>EU��H%!��"D/G���a$�F�>W��:n��3���^L+���O��T9bX���-��M�������
�n&˽�N N��[�)�Byw]���]CD��Qrr�f 
��"6�yh�W)2����W��X
��*�\��H��HEb�"x�֑	g_��:غ��db;E��Tٸ����լ�RL�\r;U<Eyǩ�H�۫	s)>���
q��u?c���£K�wQ׺ep�oA�~�PHi_�+�	A��g�В��/^*�;�=�������)ذ�z]F����i���4�����-͐ち&���;�����}��}iن�$���B�*����-���> ��8shm��{W"v�������f��$]���@RSY：9n��
x+�0���������{
���e�<B�J�+׫������r�dY���yYK	��٠q�xD�qf�q/*2k���u'������߃���'%��U�����^���A�������JK�ey��Q합��Cׄ;��_���s�$[	
��v��
ZURK�o=���µ�2~I��p�x�f��Z&%����G�P-em7�(EE�Ec��^2�C��䙋�096��y��k�wT8hQj���_�22-�ZjP�l���.�����bKN���G��h�X�ar�i�[|Y޾iR�#�Z6��.�u�z�r8��P�ˆ�U�3�sZ������te�ID��u��9�)�n��/�KRBYLc����+�4����v@|vK��Z���#$��5DA?�\���0 �TaP��*�S�ܵk�����̬n}ж{wm�ol�|(hq*MU�K-p�?�F�WWϠF�9tM`Ж��G.3�F ~��4���E�3��QZ`)`��~��*)����8n�7R�|N�
�AK��o3L�{���XJ�g �j�h��SY�y�6��󌆎��^�Y�!��7Y�?sꝕ'�j�r	p�9&ͨ# ���e�F?��QaU�w9�:�lo��ُ�+oH����+HYN4��J��w	�����*��t�Ͳ����:�->^��2(W�I��cQ`�8?*r\R�3�a��B}����JZ $jKJ�٪���A�G��7�)�H!�]xT&P����G��������k,��D���/� 9�`�}F6�|�}|��]y)/k����pD׆��՛�0$cE��w�I�bQ5W��3 �Z�G@���Y���#�y�<�o���%@��p����w~ʓ�[���M1y2�J,>�IŚ�4�㦽^l���.��]��~����بW�5/���:z=-������pq��b�I_�;b����@�,�c���>d�5A�y�8�͍� S��vlk�x��ȿ!�S�Kw�3����D`�	o�B�X(l�G�b��:��H
[��"���/,Or�/nG��%��&C�m@w�������u�f^���л��?0�ܾ=�DF�刽�y�>�&�����+��S.
�	�W��~��Vw�/��ǜ��,�OQ�房QF=R�gD��OƝ)^�-J}��m����t��8f�HR��v���(��wVj@3��/EQV�Ot�?�T	�����V1�[�z3�g�65��Nig�!~w2�aQ�^,�hDq��,_�<���ן�&�n�,�T��s���Y��NE��i�Ff$�c�"=�����*5,�)��y��O�dߺ�����:�(p�����[���T|rͣ�/�AOە`?�P(F:��T�W��ʧ��t�c�ґ���v�]5F�n�l��W��B������{;��t����wy��J���c&���i�`����{E+��PQt�S��S��ʻ'�\���ڄ�@T���P�]XL�\;��!pT@yU]�	�+�����IZ�rʥ��}{��إl��+�*Hѱ�e��0�E,��#��Rx���N=n���[ep5���mVuR1c��ׯDm!��g��e���Ⱥ����O��т~�+��n�L�Y�Hf'�M�Z22���[@��U@��h_�x1ZWtU	�����;��H��Ͳ�O9�)/� ��
���$� � }��|�R�Jh9�'L�N��M�RyH?/	�4n�d�;�0�>*���w�]/sq@TA7�~-lq���I��������--�9m�gΨ���@g������8\���w.�M'f˦��2����I����ߕd��,ܯ��[U�x���2f����$��xo�޶{�C��zD\�Z�s��r��� ΅�_�c	anñI���7c^��.�L�G^�y��u����I�
~`�/dRJZ?�y�ɮy���|�Oo��!N_�50\��lO1����m���EK����,��>�5I; ��#�A ��Q�"�m\]��u^I�B�ZB���Ý�X�]3�-sL�<4L��uYH�h)ͯ�q�5�y�]"�GΊ��݊N��K*F���� �q�#�+����bC*�}C���q����N��_��yY�$r��@��y.E���
/,����Ȅʢ�燒S��[K�����!�u^�5�G@F�/��ͺG��W�w&���������>����P���3D�7j��k�Z�2����Mr#gi���i���^�,j�սD� y_�͛��&��g����q�E�R�@b��n����x�T?�Rg�#7J��:&_'5x�n�l�e�w�\-������'+��Ej�:pN��FbM$³@��a�,�����z�f[�b�:3C��>�`�Jk�:��E������d,�?����D#�>��	��g����<���Ї.�]���gHzx9���C��hߥ��	_1�[層��4P�aΖ�펏�ݚ{l�R�c�tB����t>H�j`!�h��c�K���S7�z�g�"����)�t��VB�;�(��Pjȫ#@A@t:%�05�-��~���!�-�E˟"8��!�2O��!@����8����u	D �Qr {<0L[�$�{t3
#�{���ѳ9�-�6��ݦ����G����Y_�odp	T��yd��\�]�l5�zVש�;��8��z�I!J�.����N�=�Gu�c��Ű�#e��/�
K:�l�Z��Q`�c���$e�F<���{w�#�M�p�>���l�&����m�w�x��
(Q�
��A�h���7�3G�#ʬ�a�M<7�ܑ�~{B�5[Ǩ�_=0�+�oP�ѻ{����lj#�5��#��`p���f�ժ��x_����z�?&0��-���J����F���]bI�V��}	y���
�|�qBC��5� ��Q;��7�����*��X����b���&��I	��B��U`���hz����r�� ��@$���ȁ���A��ge�����;�[h��-�t҅����ow�c!�⑧}�[��<��g�]%`R�cK����.0:��CǾ���@	"��g-��p�oUZBD#.u2�QU���V�4�Xٴ�tt|�p�^M�֭�h�TZ��o�G��Y�j@���B���Pg4�5��x��}��]����l��v'�h=r�Cte�@�}d�;��L2;<f��HX�m�`������)��� fi��Ģ��;p���a��[3����hQ�X���jY�Tvxp1���Jų��Ua pn�x��nPT�|-$�rT<�����RI`U�Ԃ��`Fy2��E��0�H�����9�zJ���p�.E+��g�z�����'�?�R�qk�m��zl�Ko8�C���m2�VW�bݴ�$\'h�̣L�����I���CB��*��3�8�v�	ui,�8�j�f�A0�$����|ET�l��'/'[�v6�)H0�x�,��	}��j���{#a��q���z� !C2ktPо��u�z��3E]�$ڊC�%���Nֱ9�m���L���+ή2j�&kTܹ�➰�X�pe�%@����@~��h�)�K�V���I�[�s2�D�g��R�>�cA��1�@9;�I"�M���eQz��F8�@�	�'d�vҏsܴ��	�M.ׇO��I_sΏ	�=x�֨D�5�Je2z	���:dW/�P�M�g���kI�ü$'(�F{-���X�K('��EI�/��!�ڍgw`:"���CO����m����3{�,����nL�`�%��b9&e���w3��S)�{cV#�)���c�A��
 &qk�՗�W���|븉��1RC��i�� O1�<Ԏ'U��6�5u�X�ڨ�O0�WC 
SR��!+n���dT�@ҞBU#Q�*�6X���6���a3�$"�R�k
� q��+����QD�֚ L!W�?zWOM8��l�N��i9�V%�ps���17�dA�C�sm�&ݠ����]���¬:QM_�ե�J��	�-s�{����y�ɖw�|�ym�3	�tQ7���¦�
ƞ��8;�?��l��a+����SQ����꒸ 1'�k����0���u��uX8T�J A��r�`6��ݣ��k����M���t�Oz�r�vdH>f�SX�3�	'��/G�]�h�sd"� �9�W#3d��NL���)t>��9Z�1�)y��R�=f��7���r��,��al��Us��	��F���o�� �_���/ϟsE����>ғ��{�P=W�|�0�ċ�̢<�&��w�儌���6~�E,����H5����H�/�Ļؕ�E�
P�ٺ��F�8�E�)m��?���Փ�u<o���2RSiD���3��]2a�m�����T�����U�W�+�!Ф�1^SY�����Hm<�e"|��c�+�o��>��-GG�'�Ǔc��W�L*�J�ƅ�_� ��1�^q+�}t�*�.9���E�w�S��4Z��b��{~��(@,5�aS��Ԋ��!+8����:�<�9�V��8m�Am���P6��c��Ӎ��Kf�NW���`X��R�EԹ���e����/IGB�B}\��w��'���9*�X�b����(�3��x�yC����5���_��� o�'�4r��ZR�}�.J�7j�7�8��z����{����Y�S:�#?���T6�y�n��P�LH@֊����[9Щ���6[]�1��w�#_y2�E�6�\w΀h�d�z��'�h��ㄦ�g[��wΓ�}]M�.�T<��ɯ]���$�Lv_C�����kC\cmy��K'	y�\�gY�֜Uy��EIu8}�][���g�
b�F����##;�F�u�vB�������%��a�'V��Z�|2q5E�m��R�{B�
k���^��H|P2v)�H�T���t��F�_��I�@���9wЌ_2� �z�r�b�T6;[��
�b�Se~��C.������G��3�I}$����-{�l"0=�e=�P�+�g�
�������bHjYːݹ�Q�7��6�$��J�I2\��<h�~�ս��Elsfڣ�t���l�f �^RN��&���s��Kk��E] �~{�7���b��
->��k1ծ��%;U�x���L�yz�g�\Ӝ��4��Xi�Ѵ��B�2�aK����xz��t3��b����c{S�-��jP$���q�q/w�I��hX����ded`�����Q�0�ze����7T���keW��J���?y��3-6�dM�D�f��L�}���Q����8p����B�;���i�%e-�� l�$��i%�
�{�wȵ�%����V3nS�P\Tj��kL�MβK�:_��y��9��&�V�z�m~����G˅�����oL���EܥuTF�`����<j{�z^�Ո���K�?���,,�;iE+������S'�E_�n��m�^6�pơ��pJ�}GV�����E!��SA�	�۳��b)����\a�ID~�{Y�F�؇��ٹwo��cl�ew;CY���S2�x�Ѹ�-A
 �;o�LZL}�}�x����.�Bx�����$��������?���		u+��v��y`�c�Y �{�	�q�n~ՠ-0��l�\&|�q��b˄��q��9+���UUhZk��� ��54���&_��知�����c�;Q�N�ǿ��-ǔV��~����)���<t����SxC$��4~��w���r�����&9���� [�H�|S��&Aq�d��,�Ǩ�j=�Ο;&y[�xM�P�� �ɬ���'����Zζ�q��4fyM��b3����JK5S�i�U�U�0x�Q�{�8��4"�����S�q��"��r�h٠����x�#��i~[�o��T��.��"]���|�CM�HZ�<�D�Us�-
�7�RވV�����E�/CtG�I����x�	�dU>sMʸ�9%$57�a�]�Nq�ђ?�
����%���2I���#�C3Qm!�;��"k�~���p:�`:�{.�"`u��D� R6��å��ꊻ���L���M����N�2:s���Tߛ�B(�����;��UB���=�6�9

/�Sѫ�M���J��?e1���˲wk��V��/��}5��e^�����v�\���C�cN� ��(,b��q����ʩV'�֭�f�E�Ww;j���Y�K��?I����:hNP+@�f[4���u�B�qL��?�erE)�&ow���y��2�g��q��.��|Q�$�ͨq��k����¾	/а��p�Q��i�3�4����+��aG�J���	�b!?�t�{e�_ٔ�/�T>�R��?�W&t讨�G��K�0��֕�ԒNm#�@�(��a�Z[�װ��JS6���H��&�L<���pN��97ںݘ�B��d��M{h����u�7��/G6�K���fQ����J��%�Vb�c��]7)�"�<&�����]�p����G�z!�s(H��t	}�}U�c�s�@F֊�׳�'�2�d�R��0��*8�lX?u]��@�Beغ�}��c`3�x�^���'�	�"���};���,ds�k�U�5g��͓�
~b`1�:��O��w;���J��ݯ��3����Г$ˀ��w=�ROC��G�Tܙ3.��A�V����'��QѶo��QГ�s�i�M3��Aj5'��'�'O���k@i����VB�%3��ԇ]i���T�+�M-)��q=�Ƣ�B�l���m~��ҌQ�t笂�%䬬4s�"t���M�b�[+?ks���g�$(�
�����txi�}�"k,��!�9	��9lN����e�� /�,�I�X2�"�����B�g�w�wNd%���h9<#?0~�(�����)6�#�_슦2ex�"��yO�}�&�C��D `��@�S���32Qt+@v���J����_eq�+�B�
W�P�m�,��s�n鵝�V�cX�����@�s녹�z��k��u�n��Q����M?br��^?��yݗ4����S���F���4��^�Y S�:{I"T}[&���o�^�i������i#�'jl�~zۙ�QX_'
PEE�N�(���߈}����+�����|O�s$7��*��x��� 8��Y�"<�*�挕�CO��_gndQ(���o�����K�-���ۚy��-�bA��D���S�����*��}	-�A�����܉S�����w���8�"�D8�(�v ��#�bj9B���nF�_�5`g��NF27�{sFa��c[Ww��	�(1=0��t�wjR^��$��{r�%w�io�=<s�����Y�#����fbz��g���Y�;��cdpⓕ�nb����
�su�6 q�Ą%]I����o��H3�ԭU�
h��O:��i��tJr1L�t�6���Dm�.�l�3��y�!arB�"B��c��k��B_���e���Z�]��hf��2'��"�h�: ��AFKq�G��H��h4ˆb�tS��g3��;����X 5w�zx�Aۻ�6}�*�B��O8�N���Rr{8f�7����k��%j��i�nc1͹���%ێ��mC���� ~�
?�x�=u��G k(��6����/av��Z�p��f�e0�DsU���N�(q�5Fb��� HU{��5'�;,��M�p-W��D _�$�N�U;�;�x�Y�2��i�����۫{����������n���gg�g�����ž�$ I�AT�we2e�;J���>F�%YE���ٜ����x�����a.�r�k��R�Hy�o�5�om|�(��D<|��0ӄ���X=�
�.KOK~F�č��'No����kl��v^����3��9c ���\%]K�����@]� {"_��3/�)`�m�;��2GF�A:��ѫ���K�$ݷ���ήhu�S����f��% �-��&A�c9PK��"�Uf�C$��gf-n���+�ń�$��֏��Vy�)x�.�m�� A��bݝk���56hfh��;�]2q��^>XL�B���,��{ �ﺲ�H���/-�׌k,��z�4ZF�7cO"��p]r&_��J�j��y��`�z���h��Vɠu��z�����@���"<�x_C��������m���wh���O���������?��ݙ��n�����m|�� �`0:Π��g_�+G��ҙ0͚X;Ȗ�a!Q�䂮������K�'x��@А����q溰��q��@?�X�ga�O�[ӓK�.[fcW��'�إjާs�a@�������S�g�$�yJ�_�p���v�� 0H����3{Hj8�������������ˌ�~٬RL=���P�����5��7k��0$�c�bR�l�Ͳ/�u����K��;p�Y�`LP�M�z����q�L�ʈ�"�YQY!$�t���d
�x8&�$1�>dp�u������9ʰs5���W-8'��^���}�|(�U�����C|�Ie�5�F�?�O���͈'BZ��Sn1fJ�s�+�vQ��*/0�bYW�{U>Be8��_�����O�qH� ��� m7�[	1.+%��%�d &>�O�vǀ������"�(��wf�qx4^���K��A�k�RFm�&j�P���Y�p;�U��(�F��Ǎ��G�ۤ/��v����-i�E痪'�k,�6������u5�rE���&c��Yđ�1�݀�����l#yi�6R֊��k�#4��(>.�n���_	ee2���������u� �!�������Dt�זߡ�m�~7~4��!��?����!<5�Ba�W���Er5$����LRh�M��I�L�Y�uvP�|8�#�W>�Ve��wV�0��`�C���ڐ&��sq:X)���]N"�QA�ŋ<R�,�&��t9�;$�~ӌbʄ�
��	��p��n"�|���z��"�1�y{�������K� # 8-$��_}��(��z/�/jk�QG��Fߡ��\��c=����%���z�z׼8�Ö��4J� �Jv�ɼ��UfJ$
��Y���.�-��) ͵��V���\-����Yj]Mn�e��b��$� ��x0XKN�)��:�vT�z���'l�K�u�,���K�� v%hAG6�����K< J{�M0T��5��?1z��%�VG:�ڂ�4�GT?�^L����<K�4�{����u��)��4��H�g���C�v��G�2L2�}6u�5�Л\�rqM�C�g4�yQn�o��w2ooJ�-�L҇�ܧ�-�LÃj{�M}����r2�Y%N	�]G�����T#8
�JTHƍ��@��8�$]S��;�+�8h6�X�r�fG&w����-n�~�kk�er�aB��3�'>?eN�a�#Ї��o��b'D�M�=�kk���v�@hyB��,=�	��?S��"n���J�_��o��<��4j�����\!�X�����\�!����+aU�7o&�z�@S�\�T���X[�tVku8�N�n����>t���4�
�����q-����F��Լ�!�P嫳9�E�5[�O�4��F��LgP��Y_Z��쥅���N[���8n&�:a�$����(/{�#�������"Ӌ�ۘ#��F3�9�MFʣ�$nHV�Q��'�Ӟ8ub��o����Ρ��K�����j��敛�����q3��L,�شD�p�o8�����~�ɾݹ/DG�[}H��C����7vKvE���՞��>��C�`�Lxߤ)�J�t����I��Pͭ�t��{v�B�s@��7��C+�C}0Ӵ"��.R���)�XOJ'(Xp��M�VS���o�\�d�椬��R��7�1��|�6Z�P�)�� -������ǌ�/�*���Pf�~�����ęNhi���2��B�5ll$�9�wNx�]���о�����4�R�󛂙_�\�m3M�0���~/��&g��C}�e�������z}ľ�L:\c�/�^˥IJd��40$��C�佯�޺�-	4D@�������}8�ˬ�}��ʷ�`˖����s����� �'�/Ƭ=�����Q�����P�ٍ�Tw��O����z�k�w�{i�ˊOdU�l��9$%������ sm����eT�1s:�a�h�u������8{��f���Z�\<@|�=�%���f��8�YҲ�}���{�]f��Q�
���69Z�`��/Dy���SM��R3���IU߮ڌ^�C�	�wֻQC���KUh��q3�	���h����CǠ���
-4!J��?'�{sHy<��(:rk0U9�ח2YH+�{�	��q�U��c�y�b�4ˣJN��s˒K|sd#:ZJ���qj�������&�'�F�O)uƐ�id@�*#T�1>l��zZd$�mt�I���{��Ω��:���J�l�	�eD�l�(�G_Xg��m�zY=��� 㔊FyQk�̂��8T�a�;V��D�I�$FƩ�0ȡ��Yl���6���>�?
�W\�~��5�6yY�e���w;����M\�I��D�V������95�'��>���� 29_�^8��4R�oF�a���2�f�t�+ d���Wt��'ͺ���H�񷀘7�+�k�.' ��`���=Ӝ �5+}6/�_���u��3~�-���W���Z�Տ�	� Ì�u��Ml�����/���九Qbe���W(���龕S�I�f�eu<���{��l���2=/�ً!K8,�E��B7�¹�w��VǬړ� ��ߘ�U�
ۋޥ��ݫ�n�L�<P�8^�o���W7'�#�]���,`��|x��F�ɣ���n�N3�����ɩ�:[b57��s���naM�����H	�`��c��C�]E,廔q+Լe���}�߲�Pu����\��<��0���[�/Y&�iu:����I�s��x�|�x`�6Kx�qG�H8N�l�>d!�9�j�=C��U���������j�GѦae�}q9��D&�b�N���p|���2���Zd��!0t���m��ݎ�<d��9ؙ�M���o�5_�[�GN��/���1\��7	l�y��J���Q�[*F�b����
�L�������oH3���fo9�o�b�� ���*ii��8"�t@�M���L^����A4�4,
 �ҭtG�W���_�&�u�Q?R�b�Y� o2�'`�^_Z���%׵T���Z�� ���.�ka��4�O<	�ܭ��X�L6�<� =��X���ҋf�]�e���)^��lȬW@=V^!s�P��_|7�t|y�>�Al�e�jY<*�q�vp�e)t����qD�C*Ԃ�ޜ�v	���k�_��{��=�L��@6�s��W�Hm�e$��^G�Ed�2p;T�<�Vw�`�Xr���
�>�E���bs���]7�pˈGU��t-��L�k��z�y��M/0	D8>b���{�Bژ6��k�*���GAEt&2�^�W�g8I�z2^��>��E�"6�
�����6N�he���Y�qY�d��?r�M�/��p1��b��6�6Kb\	�:1Q�{����U�5�B] ��@�p�E�r�V��)�l�4�q(���<��f�Kn�����Y�(\�oXP�z�;>�*8�#��K�p_N@,3�n�9j=V�R�"�7��T�r�"�B=���Q���B~���o* ��=�!tcħ���+-�P��^��!�]��%�f�o����cb�\,��\����v�I�`P�_��Σ�cF�W9���:�DM��lmA��Hⵤ*���(����[�K�Pi@n�	={䏇F�U���`���c���Q���]k������=-��`?Du���&����I��������Y�����J�'�
��ȯ-���23���`�4���ý�N��p��9�{�1_�s�r��ݤ	�V�|Hɯ����@�B�O����ZF�D-�B�v�r�]�l�3FPD".���J��x3Jj�,_�U��&_�A�� wE-@���(�#l�wHΣQ�]�[�4��	�r�$�D�K��@*n���PE5HmӀ�jXi;FN�Jm�z�4��0�nR�g���/��k7U�Q���s����;��(�ŠE��8s� ��q�[�Ū��(=�`��@P����Z��t����t �O�-�V'o��,_��d�Yjmo?�=>\^�^�QZ���"�`$���%�p
�70����U�(u�H�Q�ȫJE@�fFM���E2N��]�0��56)�F� ?4����E��a��y��U٩{�����O���ZO(o�gp2�c���86 �qD� � �~/���ew\Tׄ٨:͒J^�'Y��ܔ�\���!Eq�8!(ǣVD[`*��&��Tk�|�Π�f��_4k92:�=�cMhZ�WXWG,����" ��#�0m���U̸5��D�~TǕ��t��\��|i�>Z��N0��%�u���X�|P�d}�3׀������LD��Wߤ���[�@�Tv�A!��7�-�?6)��Ċ���;��y�5�S�S)*���S6��>�:��~�s�쬙Ꝡ*��l�E@k>��ev͒uC$2�O�M3@�^X�x�G�L�F����̧������'��M%��)��� ��(< �G�ÿ��5��X_Z��B�Xx�ܺ�vudOê��p��S��@��F)���<�Р�)�	q�þ�ِ��ͥ
��1�b��@�`�ͥ��@Z��e������붸��x����ln:k�3��m��4y�5-�<�S'a���pz�e���%\�~!27�v2�0>�20�)�dиse�B�v�G�H`֙uɗ�����_�!�}�
"G:��A���mEf��i'v��s�%�����d��ݡ���n]�_/5�zϮ��xlo���,���oTg��D�jI )����J&�UɄ!�9��xIWР�������u}����t�_�4K֘c��v���a���1d��ml\^f���t�1�1�L�'@��g
/VsoPAo�"֠���7.'��݉��ʕLFy2���w�!g�]襠�4�Gy�����]oh!�j)��iJ�ك�U����L�̌��%N[q;�u̇���kŶlS�O��3L+�^�X�R�&�	���~��k���Z�L��B9�F> uB��e~��`�͌��cB>���$R�R��!)Jh����6;�O��{���{@3���¡�U�l���gA��7��[@3�t� �7CD�;��
�dT��s���6��LL5��f{�@�+nN��8|�2��.H6y�1�gA�7��w�S.�v|p�"V;v\�&6~!�s�E�� ��.S��[Q�7K���~�Lb)�A!��s�\�zO*$-�[��;��Ms?�\u!��+p;��1;1gG���z������]ӈΈ�Oھ��NSZj>|��Pu���� N��Vy�����oU1'0O��(J"���M�/E��,�$�v}�+nտ������]2�v����D1�?o��X!�����p��-��d:֜� �h'Z��W�^&3�	�U�:%�S%�ukxl����d�u�ݡA�x���v�$G��`�;����Nb���,�:��A
��
�WkШQpl���6��Y���+U5��*�[1�8���3B�H
s2�`z)L_�7;���X�k�eD8%w8�O�M�EE�1b*�C��0�s[uA��; ��I�(��-��2I��r�B�����dRA�z:�)Ä�;�(͏�郹��N���w�5]]׆��c&�xg���F$[��T��*���M����qxq/�`^��� F<+�Ɯ���|�@.=*�}|��N��2��ֲخn(���Y�w^lA6`�.�����o)A�������edf̤�`�}�d�Śޟx�m3�w�ܘ �
>�<*�,�e���]t~?�!�Ӳ���^T?����v��Bg���'�a����+2�?�I�[n��s7�Zr3�ʑ]cK����B+>h&������I$��7�a�ni�T�� m�sC���;�OT�0A���vk�c����8!p�`V�I��vǯ7|��ZY���]�{�p�����܂(������M�Z�z����A�Uy�&��,�zD����Êl�gy֭���0�@���q�J�Ez��ݥ�����X�by�g��T`���b(��U���]q�;�����"�(J�ə��ь��)3ao�}g׍D}��_�(�\���GFd�t^:���n��؂�{Ƙk'�m9r�;I�r/C��28ޡ�)Q�ΐS}(��ۈ���>�ua.�֛ݜ�Ww�|)sx�n�q���Y�M��=zZn�]7��GB�]A�%�*�4$TG��ג�g�-���aމ�	��շB<
;�n�@�H
:�(�/l�1��~470�d��Ӆ��xBU,��CV�ܐ���S��H@��ܐ[������ʋ��&?��4����B�����z��%��.2*ƒ�{�>�#�Z�u�������ƞ��-F׿	r\?n�ypHά[A���Ĵm�ރ}r�`�	y�~̧c�@&2/��L�h�T�#!ޮe�[��\�)9C�w�9. ���Z�2�R��1`� W�"a{��E�H�a�N�������� �X��b����窎�m iK9�8O�U}B��:�C��Z0��q��丅���;�p<Q�=n�U��Gm_�k=��Vw{W<YJ�T���-��k|H��Qȼ�-W��{S!<FXO�d~�E�Y���}�J��ħ>�_���*\��gx���c�S��� ���*�ܑ�0�]�4��<��$J��wG��m!�%�{�+�%�Pң���y.�V,�s��0pn�J~�q��r���{du�-k7�Ƀ,�<��4�)���B�s����ͼQ��%NO7��	y�kq�P�8���z�
ZD��Ia��E:w	>9H'��l(��/� �07d\"�Me�U�~�,F\_C�rN�6F�-]��I���Χ
� K�Ӷ,�	���W}¿����G6̻'�=�����PV}�;�"d��;n�=g$'�T��5�p㟃����3�������-����N>�.?�������0w)e��1m�ײ�
B ��D�]oΰ��A����'N ����z�D���[�l�"X)e��gG)���ד�e��1�����(<(O~2{d]��3/ӹ;�������m�~�ᕀ7E����L��&����b�A:y���rD��q2˪"4���'���xݛ��T���|��B�N�%\����
��xc�;���ְ�Yv 浂��՟7��"�	�C
4lhƣϥSę��MP`�|.z���{�1���[-�Ac;�q�=��*�ruCL�/��H �a"��5B��AQ��ؐ}�j�y���9�i�N��Q�~%���px	fyT2述�����e� |��$>=���*����?�ʱ �Sh�}W��2Í�P��Eכ�g(���p�fe.����s~����-��Y[�	1��4�l���A����I;S &gJ�̢1`����3�IZ�_����8;ƃm�v.�;D�P�5n}ܑ��/��.毊#�$Q�y�@��C�e������?�s��`vQd�1�^(˯��$������
�zaN��d�\�ChԵ��ӻy�a�=M�|�`�UD���B�V��UL� [j:��.O���0��#3�R�оɪ\�I����ei�k����2�J����(xG�r��!X�n���č�O�H�>a���/����u�3uF���#+D�~�#4>&G3\�b��i�4�{}�"�����ȫt�([Lc-�,�]�%�%pjL�X&�/��y�H:#�~]��cWc���,,ji'�.����ſ�X��:cys|Q�N�j��I�_R+��Q^��w�ns%�?��9�&�T��Son��N���M�2H���4���5}�xk��d���D�O�5%�^�~��C@�'��7���s(N�9x����@jI���/��NJY�O�j�ib{A�^�^���Gҁ���*�7�H��p���1F|&��g�K���+"�&8i�~4q���S�O��ƥ�c"2'p�8)_�]����_rg^�����"�e��E�݈���~	a����y��i��݅�v}����
�?�E� /��x��� ���M�\Ϸ�9!�:i3^ݥؽ ��S�A����WN΄�䓞�T)A8��e��Ƈӌ~�q�Z��kN������A��a����z����@�����^��B�Ϻ��q��=$�py���;=��<�����27u��n}wm��� p�L(�Zj�]��6��	^ݳ�0(<�.�h��c�#C=gp��G���r=k�y���i�dK�	��y�f
d�{������@��u�U�k�č��{T�J�49㬴Gۅ�:�6�>�˒������Ѳ���0��M�ݟ�ݮ���a�;��(˭��QV�9��x�'���*��;�&\`2�)�.s2�P��e���:>Vִ �qn�f��0��p�pܻ݈Q�R�G�������9p�3��տ���'��ߑ�x[y>K6�.�"d���>H�&�3��t��
���Q(�n�� r ���'е���6ǅy~N0��|5���2:�aC�:�6Ì���2d5�Kc���~�J$jb�5)�	!`�@��|Ҙ�� ��DbH�dc&��T��+���4Z=�nԙ��m����wY���c2&��U�¤r�Y�}�oT��z!4�B�5׍�F���,ۄ�t������؞ba
�oj]���=����R�^��Ͳ�t.!$��_AT�MW[�%�v�C��6����iSA*��C���=�(�d�"˲4?�>��_(OV��&����Wd�T1��mk �>C�.����_�_��<� 	�)G�Yr9��\qx����Ϟ{�ґr�M�H�Tt4�R�R�;�ߦz���FN����.�)�\�Np�i�r�}T�·�f*p�s��Y�/k�r4��VI� !��*Lg���tm��]b��p0�(�#Cz�0��w��Zd��
8�Wj�$�ZՕ�<j�D݁�h�8��y9�����A§"�Ԛ|An�")��
"t���ϑp?n!���`w��d��I��8�oci���5���h�H�>~����K�C�C&3:w�`VNSI���r��@��p>L�Q��?�@VZWl�ழP�9Vc���v9�c�Al�8'[��X�\�w��}��r�3 N������ ���[��^�+I�v��c-p6!J�#=��a��L�K>��~�E��o�i2$�ҰH��:jIC~{T�S�vRp�{o�2+3�,&�s�ĊYUE
�?��d0獅%���/�T�{�s����S���Yw.3�ǹ�3��#7��/EN��f2&��(H\u����t$]��}�R�8E���B�񾬆�N�)L{�zf����)����X9�)�}���p�ZJK�h���i��~(�k�R[�07�����x�hC$k����,wO���A��Ĩ��9NN�t��-Y/�z3�ȸ�6!�$iI�B߾�G�g^��3�)I��@:wY��@�W~V��;�mW)\�MaC�zP|,{��_���G|���G��{}fDjy��u=� �,��_T]pmw��JR:��0�T�[6����;�(}�jW��(�智j�#�M��z$Q��*����ֵLFQ��wJ5�LK�����)K��d�y{�_�
��+z�v\��CGl���ϞUz���}	��РE��}�c>η�� +�yN+��? )���\{�p�!G��k���!�����=��W��L�����{�ﰘ�����@����戥��J0U?�R��8�f��w.:�9@��)/��?�dI�p#��5b�Y�
�1��I뿱+����29�p�|�G�<]�@�WIŐ��TҰ�C�~��8�f���`��:ͼ�m7-��mo���t��7f�$��3,Y��������}�a�a��E���� �ؔ�����i�8m���!�P�wH�@c��,y'�T��y�-��
w��<�+�,����1�Ђo*�(�c�3�ǆ@�O��r���z� R�lN�f�V�f�
�b�t�Q�W�ȧ/(��q.�>͞� ����m����^��"-%}Z�ʈJ�5X����D�x+��I��?:K�#��9��Q��7oH�@X��c�r.c��0��%\�-1����d�a��(��a��y��ob�!�U�s>��B��ŖHR�*�3�D��N����R��H��шJ���T�eef�;$%I��=�2e�8�7�M=-�-���M�->�����v���ˮ?}d� "<ӘilR����{�l�ӻ��Tt�uc�.|�#�_��zV1Ʀy���$I�Ԧ��@��Ro�%��#��q<��|���v�~ݿ�:��-�>�����1�8W�!�?�T{�V�iօ5]DzC�d���7ԀQ���=��9u��\�ӱ�_��H6�Hu��#=*���Ro�j8���PkȹAdy�ҧQ�j���F	;1�~.�Kda�M%�}�=%�X�����p��h�$m}U�є��u�ud�1���c]Ή̣�{qF�۾+�Y���K��ե��e܆���Қ����.�F>�D���-`g��U�a߲J�1�����ŜA�,:�YDz�/;��uQ���8�"�ޏWĵ���
�;K�`X
����x�~��Q�'� cP��%z����x��cT�}04|'�#۳��D���D#J7Yն��!2��T �RPBZz��0��!�W^�BـFQ��RP>
f���8�4_c������-���yL{���Z��1��U�r�o�E@x���ni��Y�Pp쐵2Sy��=��o����Pb�N�z?�~�PQc��]��)��OA�B��D�TLNbv�Y0������b��+�UR�(O>�5M[�1�[XD�˶j���Й=,�"LwP�_��(���9̅�P�*-���[W�	h�!r%(��c�gU������b�L0����ۘ��Ci�y�%����\�٨��Z/˲%<-������Vo b|��T���n|Oh���@4&mA52�I����;(ܢ��ė��B�4pgãw	a6z6<@�	�U��9RH�\?�3?��{�H�_��d�9��'FF����o���Z!U�k,Ą"M�����M�G2+q��Yz�G)��k�fȷS1����4��Af	��ŰI �\��i��H���99 �\�:�0=��$3ip�j�F�Q6���B��v+=�`���Zm7Tz0.��w��8����p�3i�/
� �'Gy+�-��xK�'�\�|���J�"��^W�'��2a�Sqg/p������sFU�N�!,���J��x��P�mKX*��
PX17�����n=�
��jDP���(-�j�))��f�c�X{��`;$�vң?��;�Ւ�XN��=��Z�w�8�U�z'GU�,��L8�-��)�����1�3E��d���K�L��t߆��@M������`@��
w���S��E�ٷ2P�[[��*�(S*�= y�~n4Go���0#��(q��˦Oq��$QdeP[3�ncjr1Yk�T#�������y`C�lˬ������gX��M�˸R��HHm�]L��
"��C�1���o���P�kS]F���?�j�5,z�n2�#�O��{�"�Q���4�¿�*�@(��|� x,�=��]%{!U��͚w����e&*�J�2�M<���G��Ҥ�_I��tx�H�M M�m�:{njgİ�wф�Б��\N���[����N0W�u��0W,���*����TFP̈>㧹�aHy�����ړ?�Z-kҿ:7�v�X�Ś�Ҕ~ӢW���X�`Hw��
9bc洦����"�
��g�1E��$*[��ff4�˨��P�i|&����o��"�*��j���	 �t[��;�s=�G�,h�'���d,�7�c�Ήz]�����cE,)	�nQg�������XaK��⧎�{��e�{��s�G�݄p!IL��(�tR ��N�Z"LZ�󁶐�;"r��U�B���D�X1&)������Ɨ PSo��xA�Z/!���.U�&�ھ&_�?�G6=,ul�-,z�	=��X_Ȃ#�p7%(����2���0��幘���7ʁ������yh�0��G�+�K�e�&<��H���6ui���N1pHxj�+/3�+�,}���^��(�Pn�SA�;��ɪ+�9����d-��{��Pa�������� ����O��pB�+�w�`
�B���Ob�4S'���Ϧ��D�{���h��x�<������e.�e
i�5���#c���� ���i�c���P�F�~/��� ������Ql+R��
)���hoiY
���*�_�m�`�cG�음���5VhRH�� Bk�p�@�2���7�ZH	�\@����vN�\�G�z4��2 �&D�n� �DMdM���Z �z���]�BR�'74-�b(I/k8�X���-���]���XF7L=�c�H�#Q\���û�g�3�!��D�t*8�O����<rEIV�f4�?Q�>Fe7��N�	���}�V�����{~��2��^�躁kˠ��9u)�EcQ&5���_X�D/�d	�k�����e?\�����(�&N	�r󺌍�0 p��X��B�E|:n�S\����������U�Qp٣f�����ȤQ���-�=�����Vj,%�W֜�B;�97f�9Ղ�q��r�@W{*�aN&��pp���r/'�\��`�h�#Ba��+�T�_��k{+�Fa�HR;�j��(|wҲ�z:�iK�*�d�t��ج]>þ����0��ء���=_��m���4i�O*������ �y�Y�V��84�t��R��'cD4b�Fטr���$�+�CH�N�>�ܿ���|5U�}������>�����d��l&�p炛;ɨ_M��]��~�N��m��Ԍ�h�T ���ҿs�-�h�$�G���jr�p�����J�S���Ӯ[I�c�/@�Lc�[9Sa}$xu̎2M7�ND
m��hF�(V�$iY�)�v�R'Z.��)�9�gZ���?�V=�!�����5�^
��:O}	tF�/�2]�ꕪW��CU��B	�U,K��0�_˞��Y�:O{wǧ
��_)�3T<�zO(fX��c�zL�?�3D���0��`�CX�52uM��jH�W��� ��m"[4jk�!.�U���A��|(b%L�ؗ�Y���G��"��|�+kF̷����6�8��I��_�6���jF�ҹUr���C��֤U��h4�����^U2�K�S�e�(��
��ky���E�/���v�y�OJ7^^�a��5�qD�ד�R���!���{�Wu����բ�`XJ��N$�?�}���O����S&�����q���X#��bqb��̣��e��t���i��J�M\�q�Ft�'j���5F���#¸�N�~B`�"a���K<�˪�h�F�z/N�$����M�u�`Ck��G\^3�k�����EW���q���HCH6k����И�<R�Obi�P���4=:����*�x](���$�w+Mp�aK�ʴ�g�V�=�|g��g�������ǻ2CbT��v�%��4�$6K�7����[O��w����S���}`��}�*N0��O���!{�������Q�sS����ɵ�ҫ���7��9�%�4.t�0��1ڤ>��f��45e��`�N͒ 3~��Ł���uZ�.gp�m`K��P��tX�84Z�����qV�����FX��	�#��C�x �^�E�- C��>u�ywlwR��E����d�O��e��OvTVw ch!+�?�ҙ/X�m�X3�3��[_"���S��U-��uǮ	au2��e��I;���+4{a��t��$<����3�ң�k��Wu;�_Ǌ��n�c��|���΢g�^؆~��X����� ����S�������d
�7>��>	��zę;�'RO[5Ret>�[K�71_'\�8��I*}���G65�c����ٞ�+މ �2�΅D�ف�M��sÓ���UT��e�o�]�j�]���
���3�ǃ��p���J}����Q�U=�z�]u�gv)f!1W��mڶ~�r��շ��m�:��>���Y.+ϝi�CP4��1��.㇍Q�&(?��B�o2��Eب����/�æ� P��4P9��wJ����d��s����/9��i�?��6�CN���*}�Z��ۧW���_�䯠R���`�k�5r�qZ�/��x�� �¾
i�ů]�Cz�QX}iIGqic�7��Utb�2�R&��M��	��+QB��|[:����p������f���=D�yD6��p�A�þ��Z�o��h�]u��iV�ܭ���zb}H�(��d��.Ƒ~@�0n+�]Z
*����S4.����'N�q8�x���?���xv|��K��.���q��R�șiK����%B�Dk#����`U��h�̬�L���T2(� �������OL[�'�+ݻ+a�k=�C��i�m�=��C!�<	/
���/��3>����/�=kH���N��F��J��m�!�?B�V^a#�h��f��I3S�lbtd)��u�<��l�L���#�a����-�:x8���#Lѡ�il�9~�*(T��f ��rj��蘧��ڗҖ�[녒6�"�����d���@
��F�IYxy ����,2�3��4��(�
&Ó��1�ٚ���$"Q��nsbncm�S���{�@���ȑ. c��4H��&�G0��K�[>E^��|^k�9}�c��#:�d�0�*s=f*�e+(��z��?W�7�����N6�ʛ8��k�{���T�)]w�	�GN�E�c������eX��2:���~�ؓ�N�w���JN^��3N�.�f��2�5�[�{<R���}�L������o6x�~���0���Iz���?�1+��lJ'z���Ȳ�!ޯ��!K���\�C��
���Y��'S����!��L�ߋ�������_h�ź�M�]�cQ@nln��1�ʰ��G��x�A����t�|A-ɗE���)';D
���*M�8R}�^�FgQuГ�1��ĭ��5o�����Y��L��ש�t<8�AO�T�sR�!Y^w���`�=�1���}�0�a-	���*o'��*s���[�S���H,��ݽ�;�Fr����$[�F�$:�O%���&���)t��`���o���;Gl>TAg%�Ȳ�"��M�/�D��R�r	M�c�5���� #��C,��&��׍���~�v�1Z�;�[`u�I�,��=�����H~�!�=ӧ~#鼐>l0Jӽ�+����@V`l��%ێV[�8i�$Z�'�3��x'�+�.���v�����ȱo�E�oM�|�!�E�������n*���%��=�x�DyL���{ީc�^R�NA���;�����ڢ'��:�.����aK�h�*�b��DJ%K��c��C�J��)ڲƕ�22�P��7�Ϫ�^?)���nk��x6V����)ۯ����;ĵ�Fp���ω�I*�Fk<�)N�}�@�R;�g�{-֑0��]9��X%��X��C�rqe�<�ϕ�C�1"�{��@9�ł^��T����!u�D��t����sw�;^_���&��#24�?���rau[�d<�q�W�����e�t�:�dZ���V8`��)�se>p�W�6"3�9=�x�4�T���p7�1h�|;��Phg:�}=���(^�mc�<�g�n@����(��Ug�y��>G���%0K{c��Zϧ����"7jJ�	�ޞD;������-������b��[V�ܨ=�$&�L9��m�÷�u�r��Sz�sW��6h�'H�2�kM9=���b�1�P�$;򰎐�V�n��l�3)�.hǪ����t�&&2�=�$��9���)�Q��x��w]�}M�%:�
w���,�VS%���$˴*һs���\z�Y��f<�
Yo�Խ������[�s��3�:'��N90:�����T @���&a�B೼�Ɉ@DO�>��H��7]x��2�+ H��ҩ\:ŕ迬�q�j���DU<M��HR�a�@@@���5��1=<����F\��	�m,%mN0!�o}�����P�C?"�xu���f�Y*��+�6>�(�D<G��n;{�N�X�)��8"�=�%LyM�]���H�,�s*�2C)]1Rb���z'���5!Wџ�EMx�C�㵹3����=zh�� �G�oC��_?w%s9��K��@�ȏ+�S�O����^l/�ȪǍf!Wtb<h]��e�2�^�A0�s��92Ekew^�Dm��bw*�� ��.�.�,='�wp~�x��ؿ�*RLV���ƿ�I���M���W�<��H�����!*O�ƝBnmaB�R��r��N���/*#yt@='�j;��`ſ��D�v�90�܆�62-�R�ac��ӝd�θ�n����@�wC �dm'f�dH�]�ėw1ො8�� �c&U�>�T2�efh��β?��u�4�2u@����t����x��q��sv�rn�
6�J��$WЭ}6m˙Ja��|҈:A)E �h;�o�����Z;�`�6T��p� �H50Zi´��0*����z����F���DǱ��~�Q�2��X�V�Ѯ��^Y�3�j �%p�����0��$��
et��،O�XѡRDk�UU��p����\�9Ō��:��⺿�����K�^�wMܥ��/�f���]h�����sF���9�`�LA�?y�؍(�kG%�0��o�|\Kv{�f��)�zZ7�r@�����SN�� R0+�5~{9���0��O8V7.��G��j:��v�J'�F�ƭ�����j�ߪ^����X����P��˺���0���u��SB�3%5c�-�P�A�9ثE%�f;�a ��f�2ƬO�du���.&هi|UJ��  �W	T����ǈ ��"�]�8 �f�����d�?��ž���h]�x�D�5��X0�w����d�AKZM���Re�Xﴄ	�*�HV�|�Ƽ��*7��D~�Y�֬�,��s��S�E��[J˪�4p�2�g�v6W�P{Z<M�q<�u��s���$+�p�h{�Dt�6t���3�H��5ZI�,Fj�l���v'$�w��+k�fM)�2�O��g(��9����l�mI�:[����(�5�n�q�� �ztV�Nm�菨���I87K��ڧ&���V��Z/Ȭ4�	����@z����'\��϶C��h4
'��Lm��8����#��*���A���y�s*����|_�����!��@C��C,aU�N e�B��Գx��C������l�o��"�1�W'��x܂���	h�����
�i�dC����A"��C�iDZ�/f�Dc+��']{�;��YS�-I{�1���DXj��a)�1ק<V��]��T"j5�@��Y�����RZ�1�o�Y�9�P �:��n�f4p_,s� <4WU�-�d�4Xb!��,t�uG�ޣCa\|
s��&��G��Z��[�Mb�]M�;��7�x�yv���6�6��@ [�6>�j�*T !
�����T��:�+�ڧ6$���\�I�W���z��3�>�5E��-��N���H7����A���eGd�Ҿ��d�n���� ��bT�
���g�1�t;�d%�U& �[�~������'�+<0�9	@��F',������Y���`EKXT)a�WR��;.a�n&#��E����el��j�*w%�D���5~!�jJ��r�'n��Z\���9�Xd�e�c|஋��#|ɪ{�͟�{�3z��_���z��ۢ%�h�_}�^�%\( �<���� /�YUvSqg=-��:2��͂�`B=M2@�>�ܯX���7y�P�i��\��}z7f���΄d�*�>sR i����"������iKn� ��bA��ah�n�T���L�1��x�HU�e�n��5��V��"j��9��e39���md�\�W�q��ib7؈rM��\t8ud}��_
~����r���8��q`�Ӓ*؄U�K?�r��D��:�I�n_�~n��=\���q�'�4��k6����M�Fb|#�!�=(;7��� B�w(Կ�(t��u{�"�b�k��U��.j�� *�&�rCKY0���V���� ��5X8�� ��& �6}��i���$\α��B��t����]�1����V'�'(e]\S��t�t�V���s�Z~ǔ֭���ƏV_���)}dv,rX�.w� ������� �:+'Z�a�j �yL�{
A�QW%:�{�>�����p\��0ƞ:6p�8Io.�Hx��_����������_2a�$�Q
ae��fe]FY��������_=_��e̞,r1�E�7`����v��H(_8�<bI�fL�@����_6oS�u33&�-�u���t��Y�[���?ϋ���]���r���	��k�|�@U�Ĳ���6�Q֨�%dkW4A��xq�u�^̎!�'Ϧ�+R!�-N����7d�+�)�g�7�yU~�Y�v��*@�=�ց�1k�*_a����&��B�2��x���f�	�{^��*"+��0���o�At��(蟪��A��9) |T2��
g�ߟ��Q�h��	}�";rA��@�0�32������� �Q����
�.��PN�8�I�e�#R�糽�h_�e5S��n|�L^�9�{����j_��������F3�V���P{�ˬ�kϤМ�%�d"� ��}Ԅ�0����N���B����#}O%���%HW�0'w�kH��=�M�W���Z��
��O3���.*�bL�6�千�����N�DI�Ϡ3m�p��N�Tp��öU�$F��'���I�ck�)��cS&$n*W;*�U�s�jw�W��Q��k?����'��V>q7�>����M�My]�9ez��C@�+�RSCKnv�^�[<��
_^���O'FD���ǜ��W�u�^z�i�L��Jg�=5C��X�'Q���I,��Pd ���L�Fcԕ2�;_���`s\ 9֭�}�6@t�����c|�>��ւ��3q$]=���0�~�<w�f4�����%� ���8��[�����.�R�Ǔ�gܦ�a�cH�o�pLYw�	�H� �_��g�_P�#�Tk|�(���<��p��J�`�<�x�j2&���Ƈ6����EaIHM��t^II��sbm�	&
��%����*���� :����Bq�q�*�ރ�-�r�Vy9��� Ty��Ѻ�ݙ�b���}y �N�Am�cs��yu�������'c�6����Rͷ1?R������%bFxe�R-D^6��"��\�̙�L��̤��)�4x�e/�a�?� L����p�8tr�P�,�y<��*	��W�sV������_�G�0M�hc�"9_��d����L~t�ms=���?ĝ闷�:�,�79���P���go$9��9ʙ�n�A38�)T��L��v
x�����]2��Ӳ6vl�HW�`�B��ǲ����=O��13��$
�[~���TWS�"� ��ӓ�l�w����Ue���4B�� 8�n�P,��9�֞5�w������4��/ĜDvֲ�s�[�m� �D���"b��y��W\P��V��/��C����O���IU\8�
3'{LH�97�Ma��)�o����R�{�]�E�Cd���\d�SC�5����=ኪl��g����x��)}�H��q���>/@�?;\�T��C��a�"\K"+�lr�G�D��d(�}I�"ξ� Ʊ#��~��@�� �����4�(^DH+�f�+�X�����8�Js5ro]��ū�g��$������q��[_`y�!"����)���&��~��OC�}m,��lw�i[ͫ\w�J�E�"�� +(�`�X��Ă�v�Z���-��x1G�Ӝ"�yW����:<?����֍B���|̺ȥd&qL�n��M���/G�9*�Afڢx�eC�.��GI 9�Ob�A���-���=�ڔ�3q14� �o5H?&��n#����퇫(�~�hI��{������k�(�sc1Q &��"�`���E4;�ꆡ����Ew��|c�;2a��]Ʊ����C�OM�ܞE�F�O{@�t�ƢJG_@림�p�o��,��N���v<2� �Kx�%S�MF����v�'�x�
gο�6Ł�;H>�s=Qپ+iX4��r� �KN��E��	�S_���
fN�&��Xu�	����Us��6�6X�^W�r��7��mř"��L��G)�2YQ�0VzBB9\�'}��i��	�����������8m��Z�E4��6�`OQ߃�mu�tP*b��i����4�*��$�1�MA�S���*�]b�A�4�6�~��P��t�e��6E��F$��T�E�ZiAef�m ���2��Q�0F�g�>��|jn����E���Mo+�>�BQ?S��'�R����D���忾��]g	�$&���&L�����/�� :_�tsX�JP#b�x������� �^b�:�j�_H`Ec��{����=��x��O�����[^l� ����(I�lo3uǥޚ1._aX#��D��V���G�>�9�����%����E�/�M�oe�S x��W��t<�d���(��������V}Kќs� ����E�t~�.'��fo�p� 
#��V^ ?dw�Z�(�E<Σ�p�F�������g�t���A�8��N�r,:.�+����ڂ�}D�Nv3�i�*�3SGg�K}�[}\��Z�_�YC�R5Ql�����e��׹�D\�1!��0�+]g�E����NR���$�b|:�	��(��M{O���5� Tb���I&s\/&�ɼ��1z���.�4(��%��\$��L�c�#��Lt�Ћ��sF�f�l��w2��Cj�k+�!(/���T N$�9�ѮC�m+�	�1����G�^m��+MI���x��x�L19�"~J.>��]n�, ����1;�d�7JC��78����"a�A_˿3���D�D���� ���eK��+��w�ᱪ�ڽ�8u��f0QQ��zOZ�3��b#�4#���"��z�q����cJ)�ؗ�4P�~�c���x�q�Ժc`p%�&�I[���n������� )�`��l(��=S����Z����a/Əp�(%P��^��
_q4 7�kQ��^�z,�ٷ�t��_�Lt�ZȲ�^5��g�g��վJ�O�dE����S�u�J6���Y%�I�A�	�%{���X�tydv� ��T(,/�@G��j!�� �/\vLՃ��L�e��#����l�vn(��y�n�?mn6���8S�Dm��ܞ�>�@w���6ɨ����sf�+����v��p�����Wă�!9����Iw[���m��1E��g2�3R�������\)��ٰ�����	2�.���c�)7U��f�jf+�P�'�c��$����.�Bҁ�k��l�_��$�t�Jv�K���MDc�������o�̲BV�WX��V}�w��k!�-}�fy�Pؓ,D���|=�
�#�R�����Ӌj+����n�XTb�j��aUb�T�����s��n�i��Em�B�5:��!���oL�[ �u-��=�a<��$�.��a��}/L����p��Nݔj���V��m�!��2�-���y5Q��>5b��"��[�����4~[�HGG�(�A(/J�ػL~�oX1%O� ҥ�������[���6�$L)'�A�E�j_�x����	lqz ����M�E�HJ?���4���B��-�7�ѻ	��:rB�v�u�*�c�'��=sHlQ�W�����^"����1�j�x�k���܊;>sD���b@ß�Wn����F�`�B��a��E�Fq�ugѥcN��]��SmA��0��]Q�KK	��p/A��n�f؞��z�`�o�eB�Jiv�3�A|�49�M[�Q�Pt�,�j������ ,�!�c�����7���E��ͦ�g��c�A-5����'ե$��(���΃Tf�A�ԧ#�=���au�U�d9���mTwVH����_7(7p�&>��`3�>�"m�X�s���u�R��m�-�
����r���u�$��Xġ��c���X��k��rl�f?� ��)e�2L6�*�Q�3#�\��W�A����kst�_^ܚѴ���Xsv���zZR_a ��Eb��X�"��R�B��n�B��+����M';~I��N�\ŀ��[�<=�����
��,�7���G�A�Xb3̰��yR�-����%�O�DtIլw�T9��R��Kb�) r漗���1?��Y���A�h�[�� K�u6U1s��#[�+)������L9�<�������1�fw���IU�B�Cl� �~.K��}u���ҳHOI
���P�n��y��t,1�X���n�F$I�:�.,�x���l��?��0��1R~H-!�� �d�nW��K��Z��u�G?hG_'Kd?��