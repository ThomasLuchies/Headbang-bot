��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+�������;���ȹ�v{2� ۝ߎ#�W�ӂ����ݠ��>_g5���t͉□K2���Ec�ſ��`\_��cW��Y���NB��*�!�#-/�����0�����e	�.ZDG����g/G�lз������s�VS�]��	�_,��ܳЅ2꩙Ō��M=룯+�&HfUk�@��%��.���cm���pZ�^�&]C��l�QQ���UicM���*�qz��ZU�^u]�2�=>���J��מ�#�^Ķ���l�\*l^���F��A��N�QI�������T�xĞ��pǚ z���4��)�7�z�wcl9du�f,u���� OK���ي�H�I� ��l��.O � F�		�,& �����ͽ�`� 7�(������,\��S�!�4��ݮW���l@����1`q�f�>�U�g��E�����a�md������N���+���+���}���t�
I��-�&���I;c�C&�Q�J���5땕�?�Z|D�YP��e�|*���#܉B,��S�(����L���͙�p�&d�d�d;B�Hᨷ�ǻ��qa�+���  YEɃ��)=��������Hr߈�/G�S�>������`0&	�wu^+�#C)H�C��f�k��U�lv��v��״KOgC�Ѯx��X���8�xh��]�
�J\:�68i���Z�O	G���[s�B:�E�6M�x=	��Y�hw�946�֊0�緪&�td����q��)6��MA��PH��ÂC�&�&��R�����o쨱����.�y�l\��Ε�#��TX��j�h�>���	UK.�q�w̪V���?˱(���`�Nm ��}��Oz�t��v79W5�L���p��������{)�O��~���F3�C�Jr�)����ꅺ��U(S�h<���dk�D��Xux�M��0rG�)��)hd�a�G�{[�m�w�ɏj��Ҁ��|�̷�j��d���k�Li�����������R =)������4�`�^O�5���6���I4F!!�<�w�~��
g{D��s��P֫&��m���n��dH��B�xkZ�d��ˢ�[�Ⱦ��G�Q3���a���D��q�;��@|>{���	��jf��Ҋ^� u��,��؍��E1R�p����cG�]�\������?�+�]�Z��s{*A3�$@z�Aj'���X�0�]��_�ܗ�������ڒ���?�7�"L�6PLQ���RvT��
h�6E��^�Bz�S����o�םϛv���/�I?Y��&��;]��[�I�@ʴ���3�`�ɫj�f�T�n�o�#O�4���5�Ԗ�Vf��Gs@)ح��
��g'aӡ�U;��|X'G��O�0j�u�z�m�o��x�� =�F��Y*���|0��ϧm��j��p�
�tI+9��&
�q����e���Tr��
I/hNu��apG)�g���D�6L���M�|8h��@w~D�փ.�R�3i��U[���8NC��(�'��UЖ�^^�6(e��.�Do���j$^v;����c%����{��2�����1���	i� e�/����ӌE�+@�9�s�碴�W_T>�Z��u]�%�Y�ӗ��8������6�S*�;�o�����(M*�Dp$�&�<�Y�\�k�4٨e?���;�\i �m�>�W��쎑��!��ط�̯�f��-߹�L!��QV[�x��Ҽ�W��+����F��H�h	�����I�!l���&t*:�23LE���(��p�Bb��Q�uL�W��U(Rӭ���kӿ�Z"�T`�`�G����W0@�+l���}
P��~��qi*�h	Cj��A~<�A���lҋ�>k�����h!(��9�[MP6r�?��P9*h��F�����9ρ�2��FV�~ZV\��	e����m�8"�I���K^N���`�&�6w�j��n����Bd��L�x���h�,�Rj���"/3�\�� �.A�w�������쬑�+v�� <�Мx%���xv���]����mFr���P��}Df��Liz�
LX"^��)��܊�L�:-�ٳ�����1�	��4W�:����� �9�|��u׾�
��Mn��vr����#�~�!ޞ�B�����/u�>�n*7.S�
����b�x60���n���V�y^��8��!�d��y��!��$!����p��\���e4t��gz���|�����d�sQ�k���3x^3���M��#̌2����?�	P@�Q�,�C�S�X�jj���ȅM�ԫ�!��|n�R}��1$ff���Q���t�S!�>�� �F� ��޻����|4��l&�ȵ���1]�(8��YZ��ޘ�z�(>�{�u+{��T"���f	&��ڎ��1��~Jm�B93�iQ��Dj}_��d�73����B�g�t�����{��HDx/��{�"���:OfܳZ��P�Kf���Y���*]�� gC]"	�=A����4i�����7�^�}z�<ʉ��:$q�T3�$�[����z�h*Aw�����S�\�5�3�f��1:j�?��Z�AY-�����t���~^��+b^0_�����)��:��6��8��� zh�\����}96t/�q"�z~��w4��bNq����[��6��`?v�k{jd��6?�"5���:�Z�O�ܧ�������i�
�,���!�;Vv�$&��F@�ib��i�+�JuR�t�/�Oud�v�m��a�%����ڹ �]��Y��v����a��U��x��l|��Y�FM���{u�����l�؂F�Y�w�Qt���G��/^��D� 0ݻ	Ǻ���rW���sH��%��V*��V+�@v7]�yH�H���I�>%[ۘn� ���s����ΰi�\ �g�4'v4�9����g�����`� ��F�+vn�Kv�yLO��@I�JW�qE`���W���dlQ9����`%զ���pm��w� g�9�_�FIlb[?CF�;h�NS�`���#��g����	��S��b�Ԓ���Sk�J �y)�@k飍JL_�ג�f�p�ǩr�Q��-8�0��7�s#J@��x�]T��J�A���ϫ!d�0vxL�S3�i���g`�8�vг[�˼n�-����k�ǻ�V}.�b>|fC�a'�M�l�ѝ�j�J�TRSʺ:2�ނ�)QF��9"��F�Rmԧi*e3�}h�Tr1U�[u�"s�w�5m(.��1'a�!���v'�B�ʸ�a� |Jian!�ƍ ����<��@fdt��M�=�K*o��WX|����٫�۾�؁�2���yO��`8��_���BfM߄�uw�g�=��S[x&		FsH�6'-ؓc��UR�̦XO pN�F�Ր�%Z��Q�f UzZV��u��#�Fw�l�rp��Z�>R��tGy!�|GCg@gQk�����
��^�.Z11i��3�(^+��/�D�T��{� @޷�)�.�Z�kE��E�V�T,�ѻ�Q�(!��90'Wς���R��yC!ئJ�9�!�@�� ���#}bR�b������	O���gc�Uy�V}�`ܵ�U� �7����	 ��WBV�^),~Q���Q/�㫉��v��[�I�����=����̹�8St���
k",t{*2�A�����)w*,P٨�8�E�6b��a\�A:�q"H���G���z�َ��]Lsd�.kn�����*:G�퓠u����zB(�T�	A��P8ڃ��T���[OA1yP��\���`�W���ݷ��r�]���9��6�N�d�q$|Ȟ⩊?5��#���|��p��~���=���&�j�����*�-/%�fv$�U�^A��xK
�\��#QP��yWº��|����2y�f�ud����Y�_2M�3����r�>�r�oՏ9 )��>~�~,��\����=�?p+cty7˃O�3j��X|��&%�u/���l���H���R��s��3�;�{�˨'_"�h�E�H���񤉢E�O�r�<�׶vGږ�2��GyR%�?Ϟ9�*TPqk�(R ���o� 9Ҙ��U�~U,��?��%���7�%�w�I[r��F��T��K¸?�g�v�j�Tt��ڑ�˽��&�-��a�
f�<�B�|)+�_(�5��i���Cb���B�"s?�^�����_�+�B�JK�$��oj86ܭ��D��7%�C��n�dt����u�����Vi������B��?�a,���3��j��=e��!ۃ{�-����z���MM>aB����cLn���+ӡ&�z+Cg!������[���w���٤�%�9�X��C:@�����a��i�[��� �H!��r��s�n���B۷,v28ZF$�7�:���H(w���_�L��2�Y���CLY�VJ)ʗ��W�n�m!��'��:�{ �2�0���EH�x`�crks�����mB��%>=�g��b�������,�:���,�{������t�e�2�H&��S�������A���f/������4��q��#x�:vC�I���0�Ϸ�����)M�`
?�32�MG�P�yP��-�\�����j����핂�D�<uDb��Jr�V��%��F �����'lgS�莗��
�x��nѰ�#^c+e�d���bJ���"Q�»Q@��'%u[� �զ_gՈ���� x�@C8�X�F�\yyT���E�ՙU����ޞ�5�9ʛ �қ�����}�`n�y@<���m�;���&!g�۱�T��E����D�!cTA�0S���,�H��� ���� O��b�+�x�[!�S�;���v�+%�|?��8㷝	�`�y)�r�;ta'�6s~a[E�f��V�иhz-·Q��&��Ԫ��,��]�rtɬ��jwF�{`֞��qH	�E@���xs�㎔2]2�iV������D�rf$�d�|B�`����8Kb�"����j���vv@:e��� p��
���eD�Byd� K$�?޵	���Ɂ�(��(}�9qɳ-"��["���u��}�4e�J`劯�4{�`�l���H���ၪ:Ī~�h��d�w5���?��t�?�$x���l{��'�ȰE
:P�����G��{ѷZ�l�����b�RZ�xd�n�~��YP��e�\Ԧ�`y�.�/�0�|��|9��̗�\@H�&.���omK+c�>�c����@�ܙq	:w�p؋?��ˣ
wsB�8,�Z��c���ͨ�´p�o}�b�? ���j�b�x6�{���;��S�0853�YҜKDC��rB~@�����z��I�o��5��+�??)bW$��
jNSn<)�sR.4/7��D����D��z&�F��j55���q�zj��a�R�(�,��Z���i���e�[	���Qǜ�c5n]����E�	���2n��F�[���w��7F������tr�����R�u?��(뜓�t�
"�"�s��*�<�	��bQ}�b 5�f����KI{I�/+�y�h�D�%I��T,�N�.��u�3~B%N��_�~�%���e�S�.W2Y<a>a�	(~��#b���=ز�x-�ř<j�_����𪜿1�=ˢ�ْ��%�}�s���!N�aBF�G}Lq����R54Ӷ'�����_2������&�I=��-�<BkV1>M�Q���V[�1)�h������"�!G�^Q)Cx͂踼����:�\��T���jf0�����3����z�][�*{��,��o_s�	u���G_�'���*�_�.�$zD�(F�S@n}wQ�S\OT��t��E���k9�?؈����V�5uY��Э.K�
��M$�o^��T���A���Ks���\`���n�"^�*%t�����J�#Z�Ju3{Z]��X������7T�k]j��AW\�'�+����В|uziSt�Ytq|� ��*�AE�+�5��^��>Xߤ�5�rH��L)����T��y$r���e�`��rH�.4w�$T�P��gߩm~R�b �X2D8#�+w�=�a���gM������狟ǆ�te֞��Q��Pj���X�g�@.J�~�6xD�s�D;b�7�����J�S��u�Q��ݵ��)-�*��Ȃ,��VLZCb%�mf ���'J�) ~?�>7��#ܫg:����MSZ*2~�e���1�B�+�{Ba:�*J�Cշ�AJ�J��n�O�1����Ù���5�e
B��覒�Y�O&Cy!OE���K⵻�6�_$�Z�r�R�����V_J<���P`�1��m�񿖎W�	��L�ϡ=��� ̩�0O)���ge�j��tl�^L�Yx���WF6^�N�R�j���,O(���oӁ�c�Q�D�j�QQ��{���Gj�TH'��? �۱�]������1>ާi�nPa��&����]nd?�A��T_�ub��V��J%��K��t��:%�2�����������<M��ڵ��/\��b����q^IY�K� 7<u�k�Aؠ��6�z���u���̊[Z���
�y�" Aʫ����2y3G�ï��kK��L�m��
4�Ǳx���B�7��zU���'�H\��$�5sL���cE�b�P�T�lnY>c�P�Q�F��X��}��t��sȈz8a��Y�=&�����b��Q�4.1�

gUSV����ҷ�2�zb���a�i}QC����H{lc#F�5��-�H��@	1fIܑy�B!�}�lO7��������Ȕp�I��r����_B�XoJ�1>29g��u�Q*/�� \`�٢��L�"��d������uK��^�]��}�H����?[�*��j6`roIud��g���0�<k +��1����}��@�����} ����m� H�,�l�|5��Td�b��>��jަ8��:�Dq��P�i�O��PǾ��i;��u���e$�,��@=�n�%��e�l�ݷ��P�Jkm��sN" �Ks�[m��ee>IE�K��qϔ��Zџ~�3� ��n�̊˦��FB(�1��˃E>^_W>f�Z���&�h�>��$�!Yŷ�O����#����5����ɕxGk*�h`h�b��勸�!�!�E�U}�p�դc�2�����=��*��j�.�;��z?�C��\ �x_����5�N��e0U������;,S��yx���8�M�wB������:X��v�X�����(;���n44�:�u@� ��`���]�V�r�^\2����ǫ����c�	G�����[&��3��r�/ڻ/�iV!b�h�r�g&C#ˡ���y�4-l?�fګ�pÔ�ּ/�q�%��=K����;k�se	��g�\��D�˕���-ѓ�Ѕ�5֪��SjZO��،4�f�.���?O��4.}l����F�7���� �F "�dޏq�n��nhc��I)�}-:I�z�' p :���a���	0�xJ��9s߫sj��S���]{���E�kt<��J�Dջ������@8"iڒ���Kmc�f�cB��&ʩ��Y8[�.AvP��D�@X���yiޛYQc=�O�%Q2���m��� *�`�����)8�1��N�����"J5�F���!��A���vlG)�Ϡ�C,��~Į�q7��w�
�����R��R�^8��
�~8�= �#�J�j�/�P�C�t���Kr'W6�FS�����	��3� ����4ZRr�0h:���Y���?�ـ�^_�#s�Q�F�b1.�6�Ā_�&sD(������+���颰���%Yθ��hf�q��`[łս�$f�n��I\���FP����D%7�;,�k��?/"VD��E��.�\cs�>�Y��x��ዽ��Uc^�'�蕊�A,���=4Хn.Yɟπ�8�͸}��,��t�ȱ������rN�O'��ʋ�u��)+s�V�t|U�DS�C�V�rD�9�� �~��深Γ୒X=1	*_*
*8_���`x�E�}��2a>��Z�y�L-��{�j�dX�0f����TS2���,��V���u� ��90����h+�;�j���%��1^5h�q���BLp\1��X�S�Qt���E��B������-���T�+���G������I��A�o�[<��]�_dP})��k��m$����u�z\10�r|o��K�S��ת�3X�h�k�vS����R �@�V�<"B�z)[�_�ݸ1���49�Ҥ��&�[?�umI��o�hߦ�Fw	�A�I��BJgSE
���-��[-&��y�����&s��Z�^���������&����k�-�,'����)gg�uIu�^5*�55��<[bP�A��?�s��L#�s;u��^�����	T��	�sk<���n��{�8��p��ڜVd,���k��h�)_�i1+c4����z F)mK��C�O��>?�s�(ih5�}H����x�r�Ͳܮ?2�7h���s�	�	�|�&��Nxlf��"Rq��(��(ղ>�Fd���LG����Ȟ��s^~�I-C�ԯ�uh�\ʛV�u`W�;� �lF(!	P��=Fb�H8�����]�5�/��@�h������+��.o�	�way��Fq�fyBH)�؈��Z��]E�;��#��D'0y�g�Z����5�8
�G�H��d{! k�{�"��.J{��b�(�]�����5�g��)l�Q���}��,�'c�-�L�[X]�C�� F���M5 �:��]0�Rң�.�e���������O`�
��y ;`rA��&5>I���'���t%#t��u����byu=�';�*��6+I�X�kT"3ùsF`���v��ZQ�;�I�(ʡ\!� �膿5��g��ҕ�ۘP�z�V��l�d�,�� !�'AU6���jz8$�j�|?�e�r�
J܊'y�-&� O��ر8G���kKH�5'��������R��fW����o椮�N���#�-s�d��J)ND��W�>D��@_h,�32��9g�&_ �]�"�