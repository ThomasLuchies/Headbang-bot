��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k����W�z�N��VXi^�p���d��� ([����Um�S%��r9KO c��<>��Y=�8��2������k�h*Zd�E͌��|>�
F�1h���?���e�WNO�kk�ѹj)�Y��Q���~�x5�<uV���cBl������T�'�TV��βbB�����ĳ�(�P�8����	����g�'^+B��4��3����ki�f���M�r-�Rż�5z�S ��k(d�5WEq��G�0#�p�{�E�[��n����#Q�����
o-�KQ�j/���K��َ��"�?C���蠞�[S�ڸ����y(RI��{���� �ڎ���exf�z�is~co�A�O��&����P[�����aI���ȾR����3��|^�ϏDb�mid8,e6a�6�,j��/+̏��HL��1�(���I�AJ�n>���b��+<�!%��j�:�/��Tl�sD5�I��+gv���*�03
)����/�G���t�S���\6�`�FW]YW�Dхs?���0�] �q'e�ψ%�E��K�m3��D��D#h�+}ĄX0W���<O�Y,�3�*�[�P��*ڶ�#],�ѵ�*ʣp�IOAz3OXb�N�_4y�1�TŻ���	`t�T���a����p��_�N�������&0*�'���^��P���p�� ��7���/������|�f[a�A)�3c&�ή̽�����D��a0��S�pGq��VA��	�����4:_:��<��^����|�Pgl8SHk�1�U���@�ɏ �G�N m��R����}I`�g��W�+�Nz����e �W�WŬ���U7�w_����-�t�J_7�~�Gɳj�jz��~{�U-�Ԙ���7�H��u�ɄSXK٘���j�uX'�r����	�U�Wϧ�\�v�moޔ�y0����%Z�yK�Xw���e$�d	�����v����fI�
O��Կu�Zv�C+n+j������R�$�+(���=��R�'����G�}��$�U8���;6�$E~�����k�Csi��z�I�}h郞Z�(�ϕjW6a)�šI�$ �[�:f
���̳��E��ӣu~�����[\o�C-[����.x>1J��R���&Z]���ꗌܔ�ծ�@9Z�Rk!��d��rE�F�R�o�5ZӸ�^�g��<�"fM�X���+� E��t�q�n��>H�����J����d(�0���ٯn���M�e6z1R���+Х�����V�M�5Jo���p��܁��u�-tåR��Ƿk�G*��#�2(&dZ"�
�FUt#���"|�������Į��!�,6 6 �}EqҢ$�c��w2��=e��D���v�%,23�i�G�־dx0��.gt�.�Ⲏ��+���Qj*�����c�\!�<���{Q�;�|�!9�����=���,	��V{z���ݯ�����`��}]�ξ������tWk�U>�hh\aǜk*��_��1y3��C�[��$��c#dr���e�uV�&���7;�иܭ�9�Z�G�bF7$[��c�O�m<�;����mJ�;��m�C�a�)ф^���I�6ef��W)U].(W$� >�0<�a�]D���a8+�R�K#%m,�3�EO$����������c�����w���a�K���L@I���h?���ϋ� )ͻPdg�žm�<��Y�:�m�-��þ��s������}�R�K>N���0������k���6P��G��(sv���3~	��@1wɔdT����d�)X�5�Zˊ3�eB�py����_>��A��}����ڦ�9�Q%��?>^ww��Q�~��\�SGs�eOg=\����Zr�נ�O�����7� �GR���V�v����)�J�i�6� ڍ='��'��Q�#��3����R{��u<?�+9���G�h��_�P'i�R�2������ӏ���}����ug�\n�-�+x��G#}�;�U��kNR���&w ƦF�/jϺ/�i��/<~�t|��B�x�G&
��{�(H��g�2�-c���7{Ƙ����^6��X���񽤁��^��)]𑆏ʒp^�3j#`Y��u;s6�����*��E	~B�~�v=x*]8�t�e���|�{���g3P�ObD�g*���d�J��	�>)j
1���c�6�L�o��eZF�y�WS[��A�e	w6�<�CO�q	�X�A�?NG0D����ZZ�{���l5s�p_��v��i���L��;h�iu��m��x��p��s�����I�;Ĵ�u����́O����Ж���W`׺1`q�{����ܣG ����qn��
S1�D�YEGa)X�ԧr��a5��k���C��G�˟ŗ�����N4�-	�	��/�.�5,0�
�)���26�y�Gb�n�iF�� 傎��W/#{�׈�D����pw�Ʒ��rKT>4�$�T_<3���]:,a�X���j�Q��X;C]��_7�&���
y��y(�mqM��W�N�o(�$﹂��x����o��.Q�:p
�۾Ώ*�D|�;�S�TN��sN-�/1,T�2!3' O��<K�Fu������u�,��g{��H.a�w�Ut��)�Cd"��u\T�+��Co{�L�{t��H��}����%��Ѫ2�#�Y�`b�5ђ�X�,�B�B4w$�Gbk�'8��&Ȧ���td���n#��
l�����>���ɨ7ck��`G�v�Y��@I��3hN�5�.��������u�¯�n���=ל��\��=/��΀m�fWb��æ���	��_#W%� Z�Z�aT�z�Ё�1�%Z3����-�~�#��a�C*�+��@�x�=	D�_�[J��H��m�xA<���"�CMQ�Ͻx��M*�-�
�`��/aP*A^��㠺�����?��x䆅?�>A�3�z?�~ˉ��'�h\�j�����@z�,������ӧi�+J�Y?��$TV�y���:\�^���TV��p�֟�d%+zҌ�^`	��F`��?�l#d�vP���hG���0*2���"�7�;E>�+v����]˦یKru���>u���4G����|@.M�sV �(��U��3\K��~�Y�3o铫"�U�M��k��e]rz��ev��u��ݡ�l-E_z i���]���f��R������O������w��w\j�΂����a�]x-�P���N��9	{O%�����~������j�Z��]_m�~�����ç�9��#��@%��o7��)��4F �v��Փ���:t�n��9n��3��ĩ"��4>�۵wC7��<��^�Rެ�