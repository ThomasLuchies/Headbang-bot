��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k����W�z�N��VXi^�p���d�����3X��#�½2�Ү�/���X�Uq�UDR<�d�P��*�\��{����Wi��#e~hK��5H�"���g
�ϧS��]� 7_�]O���͔����
�2]��A/���=e�NJ���lC@Y �%r�F-ژP���~@�`��PS7�X�A~ǻ���r�DR�[!��衎hz� ē�y�5IIͯ�1�{-�0�5(\g����}�4v��?Q��I&�Dt��
�a�,|����)����b��JE�L�� �J5����9�Nf���#N%R��x��Js2ͣ~�����þ���Lu�%v��"�6ޓ�1��e��C�Mg �j&B����g<��BCy�j٣}C��<�n���q��5�gR�h�ڮ�@�E�¬�d���Vĺ�������T��!Qwe�l������	Q
��T�]�/N�[�Ǭw�t q�f{��S�C?�E-{w'c%�<&R�Oqf��� #Rx�.�.�IV铟u�8V�IH<�׬��e�KC��j04�� ^��u%`�_w�'a;a��<\8_��(p�X�Z��"و����:w�6�~�H����с��1515�wqJ���#[e�|����~�UșG��󛳢�R%��#�nrN�fg5U���]M��^��т�b��6F��g�����IpP�5���/��������K�횫m�G� ��pi}� ���C�?�r�R��;\ws������Պ�a~���=Д��ù�L�\k<����X����FIS�W}W������9��@� af]���bӟ^�@�m@�������7� -�|ò-n�{u&|:R\�۫��ݩ��$�|��[yV�c[��Fm�_o�&9��J�xe�W���yK��E+.E��5a���լ�;cQ��1���\�`,V��G�>}z�19����R�&�H��%���e����zA==���p��1���S�7��F���,�Ԝ�M���w���d�;�|�1�GF)�WSq���ҵ�0E^�� ���!?�gK��wׄ��{ޅ��)|E���K�����Ob%vK�-%��F��'�^]�|����Tw1���62$���c�j>\�N$ �W���>%�0�0��cPwG�(����hm��k7��l�K�E��
_0�]�í5�;|��5e�S��\���^A��/R����DXw}��KC�@�z4�T��6���+�}��L���MV`_�%
i2Eu	5:�~!��<}c����SJ6b�sQt��Y����4=WU	�z�;~$+�����I?�C=��[���P�Dl�@�Q��J8�@�f&�^���v��"wߜ�)F	Ϛ�D5������G��+2�/� 3.�#bdS����I����'�4lH@��f�\��,+���f���R���>,�!6��ИD<�Q�H��,��O8��7`{+�W,귖]�V�V���#��ߡgBA�ӷ ����\�Y/�ϯ��kZ�?K�{J�#�?6�����g��ߌ'��/0��:W�@z6>k�����6&��+�'K֡0k�Aِ_p�@��J����	����=d`��dX��:9_[}�<?h%�bw�����+PVh��z��m��`�4��������Z�)yhV�(vg�s��b�m�������k( �u{�Z�����H�ZB�}5_��t���*���q dO�	xl����GDH/N��[d�+r0�9��3���Z�<�`Α��S��^�\&��v�rЍ��2ޛ�_e����+2�r�LI}�i[Q�\4e6{=Xs�����ȡ�`�h�'U{S$�]:���z 	L���Tx�l��~���D���o�S=�,d�e�/�8�2������qMw��^����L��&��ML����K��=x4�8qj�w9J"M��/�B�#h�Z����20�k054f>����޻2k�d���rl�]�5�ľ@MBh]Q��(��Z���E��Mv�
@����Y� ߺhCC>�-.�`�>o�#i�E�T�8�ex	D/[��7]���V4-ؚV�-#>�j�c��_YM�7�������i&^@��ٝ��n�B�G��!o��>|�Q����}��b�fu�1��.��,⽺�i�)�L���"���Nk	�W�K��QR���`A�?-��6od�p�1ׂ��J � ���Lk9�dN<�1�ۑ ��~7��~�F�y�0x� ����Y��X�0c�r�#x�S�<yk�����L6��Z�'�b��9�^����7����D�!P!�0R�������=z�O&�ȹ�o��)�`vq�〇���Q�3�4����W�miNm�P�d�3�ϡ�၀����3h���¯*f���'���Km̐���sAH���y	��k˘h'��fF�'��1I-A��,��^M��
�՟����	����`t��F�������R]H���H���[�[���|l��9�KP�@��x���MB�r�ыsG	��"��n>�n<�s��G,��#�x�8�43ڄ����@�We�N�.HL�zO6.��u�yHz}P�K��ԧ��W���J���33��K��y���B�º��n\�x�)���υ��E�dJ)���S��gS��Lh���Ӂ����6s���>�y�Y��=ԣkm�$��7��R(�چ��I*��U���
ic��o�������C�Z��o\4�m�&G�	%`�K�ߩK�����}}�Og�N*^�/+l=������0_�j+s|���H�iUR,BY|���m�{,GB��+�$� �(t�Fm��zs�0&���N>W���ڥ�3�ɬ�낤�D$�A {:9 ?䃼�bi�Z��`��_��W����;��om8���I���53�⢬qT#������ǧw�ߋ�gs%�;*	$˔/~��Z��GTU�=ͨiҸҴ���0Bn�����͞�~f��*��`)��=Z͔X���-Ļ���������L,b{`t�V�_���I�L�Ǡ%���]8�����մ.Ԡo^U�]d�W�/�!4��>����w���(�V�R�d�7/�쑺K	�,�=6��0C�=� �jEs|}�,�>��h ��zG�9@�{����P��sL�����������b��s���ܑ%]4bR/��d\ǚ�D߃5�G�<�^�� �>e�4��f)�~K�$ &C�-�t�ؙ�\�A����x��F|��a69������&�V�>��Vݫ��~$��-�������h�� V�9ň+�$n�t�Д��g{�N[���>Z�y�Sف$����+<���&z���QU�`��.΍CLQW,P���X�X�y{bWI�C�u䣲�L/��h��Yp��� �O��F���G0��� ���!��l:�<� �4.���_��nSO@D'q�%�A<1�\�OU�ݵɜE�9�jΈ�;�a����������6�`&F�R%;y�G�=E>��L1
�ح��¦z��^(KQ�,�숗,�ɷ�M�NrN����iZ
(^	p�_q	�z�q���n�]�<�_��Qtl��.���jztiZ��Al-28k ��}QNF����d��zl[qME�mR&��#�{6�f#��4�m�F��6�N$���s/���(}����$�.�������?−17� Z��f/�i�5z�2�T�"�ٜ��~��-Z�D8B��k1�-��B�j�o�I�L-�?̈́��P��y�&b�#��:�.�n��.-
�� ݘ��2�56���@��
`.��~a>ϻ8J��"$<c���L{Q�n�U�h"�DR������-�z��]#خT�A�r �� ��*��j�Ǿ��?���bV���T�[Hm]�~T������>V�(�~_��H�A. �¦7�ו	�y��!!
*�i��>���e���ad��`��)8#_�i��N�|�tqC~��ķ�<���Sa���Siu5�]����oT�����H��;	E���z��ۓ"�kM��:H��*�:w?D]*�������Ym���VE?ňj�	��U�'�@#���~��W�윯DG�LbA���֏�9��������W�U\�;�
M�z4¨Y����i�x
=22D��Ĩ�Ƨſ��Jo_�h��T�����J����M)�G�ߟ�k���%���O�W_�Fγ�G��K����U��3s�~$N��y� �;�	�����ﷆо;sD0��������A�up�V����P�'�;�0���X`���ĝ`��d�~��� ����ɠ�z���@8d}z����˕0&ZZ��.�x�I�2�?M��(�?�}]������������p�fDp�+3�ϐ�$1��,��"f<��Q�D��a���|fTD�{��_$OS�}4-���?�%0��aD�.p�H��E=�m�l���R7/I=*�6���ȸ��	�א(2z&�+;ô���Y�r֨�����Y����n&�%���W�
�
�6���,���ʫ
Uȕ����@��͐�G�mTE�M����!��c�
�kՍF'7��{��ቂXk�_��>(R��9��Ƃ����ٟ�)�EC0�Â̳4֐ѐ���D1p�Y�pr	S
!?�&��`fbcn&�AXL�즈�O�C{4lӰ����LW�elA�mr�qȎd��1.K�_ѽ�i󦴃��n���A���@�,�OI�'foN
[wt�����zr._M7ϕ�;W�M�a�o�H��v��4������P�tS'ʚ��зؾ4�E�#��#���k`����Հо�Փ�f|q(�`W���L ��\�B�7���N�&f�Jؑj�;p��E��뜰���!kD��6����D�Q}T�"_�����x��Gu���"��Z�`�4د!9���6�8]���3�}ɏ&�X�Z:Q�m@^�� ���>am�ѵ?(@��W�s������ڰ��A����U2����#�i["3\�m~���	T��2��������H�qh��C��d�F؆���ʌ�y��5>7O#�,��j���iţYR3�c���L�j�&z�*{ z��9�\V���t}�^�5$D�p��������#����H������i�]^�9� ��K����Z�#Q���1:���Ir�����U�,}?�_���\������2�����ս��B|,�c�"��>������,#��M�27����%��n�i���ׯo�p\t
AYr���my����w�<%a����8K99
���$���@��d�c��Ⱥ2X,ƪ�,���A��
{Y����:�*�Ax��2�����v�W9#'^����\H��]�T��(�	DoJM3,��p|TTj�lk��"���&ZA�꫐�1g�KEO�\��~��N��eB����/x�ȩ��s�;oaD=ywA��@)�b���mU�㪭�&���R�X9���j�[Z�_������h�Gi�)'~��Pcӑ��AA�<�F���uD��nr�U�cp)M����}�K s����%�m�x�%�p-w��V_�͔HLB�Ū���lH �)����	n9��6��h\d��rM���M�M楽���n�Ͷ�v���Q1~����Ҧ��MT��[(r*�\��l۞{�E�Kì���V���xx�l���嬮�>�hπ��g����Ȏ0B��j�]M)䄷M���4��G�KE��*���I��*Ø��i�����h4캻��n��*�\������J;`,���)�S�,)<�Y�F�	(	�����;q��L��M�ɍlJ�Y껺�M��F[`X߭���Ge4Шp��@�a�Eȥ�c�яA`��jG�1>�L'���Ɂ�Uc��%�C�����8��3��3<��3r�ev�F+�@c�Ka~Е��7J�����8_���nĞs�n(g��p�g�~z7������0c�tFh3(}+�N,T�&3v ~����!�lڍsU�nƑ9��
�wt�ބ�:�BB�0�r��y_�|X"H�,�a�g����0P�u����*�����_�q]wh�|@ڰ-� ���p+4���Z��|Η�|
������]'���fzLO;�����B��R;6��R����*���a�ݵ��^9�����[��7��A����pѹ(��J���-Qc�����oݲG���Uȕ,�A�A�`��a�6��!�,����A�Yc,@3`{ �Ќ�g
{`?(uN۠��4�9���9(��[��(�aP��_��*z�/C&%C*q�H����ۅ����4�,R�K�l�����}�d�Y� �ق8���~�)ҔL����%��݇Կ�'�6���������ia{OY�&�s"r|�_Uc�kJ�):�[|�ߥ�q�o~��g��5��#{U/F��;J�c0�0v��m����n����`�z����w_�d���O��,=��>�0&��-V������{�O��b�&���\��AeVV��*;����%*�uZC����/��{��xf<n�F�y���f�H�ː�=���,���ef�GX��c� ��}�1�5QÿB�A�C�l��
ʋ�}�RƔffT��X�*����|����Z�L�WGi��s�Q�F�{���Ν�㈼��ϖ��Cԝ���:��"��h�o�����)
h�,��zh�b��8�y�ga����	E�y�Yp�cY&iƭ%��=šh���Y*���"u�I]'*��G���I�Clx>p��k�G��}�r�d<!���\d`� �r��_��9�g�u�{m�޹��#�����ò΢q֜����Si���Nt��?n�r�'�yH�6�����:|ׄ޷�7z\����t $�Z��4�E��R�3<�e�ZL��dp2������:l��*)'�&��#�Q�"�Et��4���epL/�����q�i�~�$J�J1����^�˰��X?��@�X�k�zm�}ڞ!Q�}���"��N�-�8��<}���F�!j���^~X���?�A�?<׹��5�BY(X�t؅�e������ � %Oж<�H�C�H����>�s	�D=�p�r<hQ�N�}�,<���ũ�ھ�;����_����*#o9�p����G�t�����mV��Y�-�i]�	����nTjKb �_ic�$�bU<�4��8�n�������?�C��"o��z����ǣ�]l��L� ��[��=�Z�t<�B�1�w�(���ϳQ>��g; �z{ p�M�7��ؼ
* ��n��?v�w��Ⳮ���6$�+��E��~LD����7�W|R�3�oc�����6�'J.~k��ݫ�c�4��R��*���%*�K��B�[����R��b4�P9Hu�o�Μ'��~�eL�q7{n
���S�@�s�jB'ۗݑ��,�qg ���"��1A�4��X���`��DGQ�T����7��S��ʈ�y�+�����vЏ9�Hע#���j��(�
5Ƌq�S0����=îG�J^�9���Bh�ͬ���h�ji�p�B��2��,�P�f�S����;��\�����/����k@=]�1�c��~�-��D��!���*��G�}�շ. V&3��W�����^\W6^;C,7���C��(yR���1�z�m��y<��7$$�5l�3'P���&]������;b��L�Y��8W�;_���5#b�Ea�WX:*)���M�
%����?� L�*�F'���QZ� ���/ s����Rt�5��t�e0��۬`�R	ü��8��mRl��\�������xS^"D�_��[<�x`�Rb[��2��|�CȅM+R��@^v��gB7K��C������\_�/f-�յ�1���m:'����^���]��>��v[�>��r<#�%�Z\TN�L}3���@=_qMQ,¤{�·F"�����xI�����v�m���dq�f�#��d �)�k�^��QAK����|�bP����	�b�du=V:�ZgxS6����8/�e!n�%^�� �r֭!^����L0}��-����\ڜ+�ʒ�H����}P�k���t��.��ϗ�� �*��!��`O�ӻ��8�!�C���4�?������4T�� Hy�9	��hc�БZf���s��۸u8١�����'V��p�25^ri�][W<$��N��\�P���ٺ����`�;DZ.��!�x�N��ҰL�\g~��^\K ̅m��F�9D�>e�$4C|r�\Ԁ�#�@�׆�6���F��r;�31;��;�k�ݲ��T%1�S�Տ���Nɘ�WR�fC�&��.�e;��s^�4�K�9���b�ӗU�f�� ���=�v|���E-�7(@�n�;3��B��)�SJ�*I�A��m'�`oZ����`�_��l��o����u Kw�����H�1�a
^Bn�9�ٌ�P$����%L��Dߎ������BX����6?��[�k�-q���rG!v/�~�����y������2��Z��T�o?6E�C��>#S�\�Z��H2�v坫��1L��_���V���XK����9��2��c樽Hb��%6�n�o�C�}���_�@X1x.V٣��=IG�=�~��>7�E�2Njd�կhd,��W�݈24�b�=�F�q���z�<�l��Frj ��`�L|��i���[�,J��l%��-뾝f���`��o�lb�T����f��>�U#�ّ�^M���[�4/Vxq��c#��@l���,��j�^��A�-x^^0��_��b�>�ю�I�n��a_��!gG|&)C촇�t<��,��F-*�$i�h҅�̰I�Ц���~=a��j�	�x�D]��fL�Z{� ��a�1_:0�\XE3�4��g��7����s�1ǅ����|&��9��V�?�G��ʔ��y�����p�_~W?�_/m�|(���y��>ߜ1����/&��#�i�n�ڼT�v�
�Ն��:�]��C��,q�N��$x~�((�S� -6�G]p�B��%:����e��VO��ɐ8`�P|�AͺJ��}l�?���8k�e��۬�Do�qI>vj ��1R�N��Rb���A�NWWU����Ϩ%��bnE�L*�րӷ&#��r�z��%O}��
"�ƙ��
p,g�	d�g
[��0t�p{�����7ݬ)��ܥZ5l͆�DE�Ts�D<JU����5~1������K9����F�*�wަ`i&���6�o���Ʌ�
�Rd�p�K� Dx�Z*���	qh�|:��8B~8�5�`u��lsǩ3�ʫvI��e~������]�C�_��D��W��i�-hi�� 7Af���qJ��*|��,�vnI2b	>_SJI���u��2�!m�	v�Vy�L��\CfB��)d��'C�$��g	]�x����|ifR|�x�0[N��J���xZ`Wl�>�{��ЕP���d6�B�(�_�� ủ��Z4x�{N�Ώߩ-���ٍ�Z�~��v}n��cy�����h������G;������l!ˑ�E��Ufʁ���2>P(:�94���]��f�rQ�IE���q�'=���?����G\q���>��l��˽�單y�5S��'���Ѡ�{7\���3]B�-�����I3>`�j��-V�˟�dhk��W���a������>u���hM��_J7`� ]�DuW���u�TZ	MF<�˶��y9w�3����(a�Dk������`�W��5*_��!�0I0���ļ�L��w�
e��lƓB��l.Q����x��������*Sg�۾��f����J3�q4��/4o;L�l|�kݨ��VY1�ݟ������T��D�`���s�T��^V^�B�VwK#��}����|�T@ޱ4�5F��8͒[y�*��ȵ:D9`��y2�NV���Db=��RkJR���$����!�1j�.������ˤ�+�\��D|D	�jY茚;}�X$.�WV�� �2�i�!]�T[kj_�2&�ᇿ:/�6V�����Ef�ڙFZ\�U|��QC���%��q%�.�r��M}�Z��� 0�c|��7�P�!$,��6S"R�5N�>��S����VH��h����$�w����%0G���/��-<���)��� ��ol�O=}��Y ���O$�LL��1���0r�Ҳ�%���p�:>�?0�7g0C�<����'r���g����g���H��JRģ��|�v����Ͳ�+��;H�>H��]���؋(�_�N��Ǝ/��l�K�4B�E�x�³A��8ک{�ϵI��Hz��w��@l,�JWE*]�F���B��cȌ�v73��(�ۯI��v�~��n�դ�A{.��a��l�B�18���L��cTOl2S6Jmwr7 ��������29�C^s�[.]�GOc�JXe7��܀�պ����m��		'�4	$�.�5�I�]�P�O
�ᣂ�dsZ�&��z��l�yn����TZU�>�ɞ��@6����V���0�����)��Zϐ?G�x�EG�5�@Q�<6�G/���X�I���j��9p��	�9�Լ��������t��l�;hON����d�MQ�O�VzK�b�.%1�����?���(-K���,�@c���O����'�悫���()Yz�Ԯ8�\7�v�����0���P��K�D��<''t���auV��ʪ���]��`̭yr9��P����-M5*��>�v�E�A9[}f���@�"!��KJ�M����̇b�	��������>��B�֘��������{�O~�g5�C��%�F���޽J�!�Ɣ�:����?;�QX+�)��m�wE��|>�`{g�o�MF��[I{�����S��L����0�󓡘O����U|.�a�(�������Vw�%��ZdJ,�U��~O��yta��G�U��̫���̀&�XǾ�4F�b+����1_�,�(�xD\<����n#�t[{�����E���:����`/�I�P�jQ��������~�~�1Ūb���5ۖ�h��4FB�\3��,M���ڊ�>�2V�4��sU%�����݁;i����7��๡�,�ַ�y������ջ8�����rp�u ��W�poe�gO�t�(��#Uz�]�p�oV�N�l�YB�Ҭ�S�D�_���_�Q�i��:�~����:�I�QAպ!#V�k5�������A{:�Fγ��o`���d�J�6D�������_����M�����k�qX�vE���-�`q�'ݪ����ط���Kl��ͤ�� �s�g$����/�STG{Hn�1�=\��v�>�-�A�&/�GꐕjL��m�?�� �9��cLȺh��G0�:��.�1�_�����=^�T
��ϝF��J?h-��E�YP�@��~:ͨp�F*�$rQ�N�lf;F˱KSx���ńl3���O�k�9�$S6O����%�m��O��u�� ���h �s
d7F�5�A�HA媋j�
��A#���c
Ű��R�ۆ�����V8�-�[���!Y����X��0/�|T*J���6��\&j����jrN9Es,���?��t�A��$�^K2Dծ�?"���O;����8���	��>TL�Y.���"��^���d(FԺ�H��ލ���1��Q�����7"�Sgu�s�"�*$Y�!9��b˷�|8I��L<�{
�LX9s��d���#�"���M�&7{�G�\�ˇ>��a r�������Ae��>��ݞ���P$�l������V�e���E1Ox�+�d����q�o}�O�w*rĲ]��6;��J/�f]jY����2 Z�T�'�2��Y�:&�G���&�wJ���CF�Ň0q���cw%KB&Y�13��0����1����D��x�SZ��[`z�Y��
1�X*���,��tt�ϥ����i�yx�?"R�/�T�y��BX<AI�+�'�)Ƙ�_"��Ƚ� �B oB�tT�6C�s<1 ۸��5@B����U�<�DxD�*����or�xI���:�<`��p屸���uB����ZUw([$�n�Vmƍx~k��u�!��j7x���.�k��&q
��S�E��$�q��/t�j|�x����e���f"�ˍ�u ���e+%	���pC�<G�R�B~:Ja=؂���?����ӹy)��Mzxμe�"��������)��Z��X��&� O5�T�Sk��k�;�a�����Q�,1�Y޳I���4h<avW�ҕ��l�H��g� t'�
�t��B��n�
��h�� �4�	s7�z�0�?� ��J������?���[�E�@2ѱ_Lɟj*#��s:��(�� ޚ���Կ���ɶQEט]O'W�LߴS��7�%|��e@r.�]L�����]����[�p��P��v}�Ө����^�1ƞ3�^z��y�������i������("	U7��a�����xu$OY���nZ~R�Z�Ē2l�O`���VA��p��
q�ۓz�N�Q�=�e�=��;��!���v��?���3�|d����I�1üL�G��y)�_�{�M%7z����=-M|���	�q�x��8aS2���$���Y� l�����ats���F�}Զp����os��*W�ј� �>����t�\!H�L��Esړ�ggCQ`�)�~��[�2:�2%Z�Sf|F#/�r%'��7��߁�Ͽ`c���\�K�Ś=���܉�mI7��h7,m��c������7d�X��1i����"t�}ߙ���m�j�=+�-�B��U�L�<���%f�W>` ��x
���]j9Yb�2KY3�}�VWV�ũ8
Z�s��4�I�P7��X�1�l�/��>���Bf�_r�EG��Zw+%�a����H����D
��~�ps�ui1E�W�H2����G�ı�,i���v��z|��+QJ*�f��o�����5LПs0���QS!����y�<��u�x����r��
QFcJF��}{�j%o���|(SmzԱo/�I��w���0G�q��j[����(�s���cUr���?�p&N��	��
z�>��F�c��;ʹ��${Λ�o֮�mՀ C��Ş�s�������d^�9de������=����M࿎h��������ǎ!����Ƞ+��>x���O���)S!�������*n;��f��Y?��G$�E�SC��^�
�$��Kl����d#���܎`®�9$��%��j|�Y�ډ�W/e鸝Y�n?�MK�c6�J�����ߡ/y7O����]����B)/���l?��e�"3ͷ3_�Ι��=���Bd�Z�0��J�V[������3������I��*끢�A��R�6���"U9K�M�^A}zO���%���zQ��L��Y�����1Fd����3ɴ����2ͪ�_�|�^����bIČ�5u_��L�y#n�^�ȋ��&��)ۚ��,�%�TզpI��l��JAK��������k;w,� r9�� �5�;Li��6�q��zV�z�%����H�La����{����^eYy����%�z3�R��@4�{�\J-���$k��v�_���R�c$Lm���t����>�{��j3��7��&Uc�'��<�9�\CO�ngtM��<;�=�����pn'5���
���VK�Z�%T�d>c���?��%8C��f܅4��TL���Ԑ
/�V܂*�Q/����0�5�lKBt[�K�tbR���p|a��H�gQ�����~M1Q@m��:���Q�$���2�A>��#���-�ћ��;7�
�:�◨�#	��R�*�r�l�l�#�|2��߈T+�����LΗz!�2h������PCt����ѧ��in�Bd6��'92�M<NO"'�j�l�J8�l+<f��sB|���eѮƑ��	d� 0����ˌ�j��8��YF�$��%�8�ވ���zǸJ��߁P���I�d��?�	O�o�?��7����b͙ԓې�s#�����2�.�\�M"负;/e/+Q�c�[6)j���"e�b-�%ϒq
��L������>�9$ a?�0�q'?ޞ�ؾ�YѷaJ�l�?��OQ(���1y�g�C��͞��mU�����=�д��
���-������V=��a7�S)z��T�_�Ea���"9Y�B���ʫcj��S���y!Mp��RC�at[�<G���rIhJ�$G��<�!	�k������!,ޅ��SQ��"S���V!Q��G�Ty;s9\Þ�]�y�&��r���4��f��$�6 �*״�)	9U���3�~aD�ɫ���Æa��˚f1Y����t�吏�w:��YU@,����/odI�e�(�-6��跸_e�A� ��4���a��P:��0�-���7|���N��M&&�ܤ��V���E'Q��@���b1�r�]��E;�W�O�-��°:�0�:�ݶoR��B�|�̖^BC��0�cny
:��G��6Z?ƹ[�:vVĝ͛+~N��#,=��%�h��$ʱ���Z�b�V������41V��T	>-�Hb[��ROM���FRu�r1����э(�BX�}ۖ�S�C�y�A��g��Z���JuD��?6��X6������7p�x]d�(TjK�8�4��ʜ㘸�?�{3anbV�A	�&>+$?1@Fbʖ���(��T�.�狿��� �Ů���$>�ߛ'�7;a�p��2/?��_Kr�"�M��<����Lo
�J�ѭ�~��;!��9��E��;!������54�-�e�\N�5��a�f�[h�
��)H�@���+rч��t�_B��*�L�i*��'`�i����E�NӤ�Iu�����nM�bi7%���Ě��E=�k3j���a��S�*x����ȫI�E9� ʤ�o�v���W'\E����3�Ɨ�!���u�����?i	#���.��x>�h�O,�3�������l����Y��/;o��朎��CH6���k���0����yU��K�����;c4�Qe3Z��e)�N�4�LӘ�������NGʔ���u�̎{t�;�ӹ�j�L�AS4a\
#s��&΋U"7&�0A��r���ı	�h���ь��v� <50�	��|�'M����K��";�.��;+�"f|�<�����)�j�9����=!ʺ�������tF�*��8Řۺ��O�M ��n��Toi�Δ�i����G
�^Ð�@u���TR���4����@eW�;��g� ���4�\qP<���-�ՙ�O��C��ٵ>��i4��l���=�^d�( D1��8��ѳ��~�5]���b�����Rӹ_�6k&��b� �C�`\҆� Z��(:���<��-���v"��)F(��N�X���n�^rzY��m�]録��WMM��Dxy���7�{��F���;�!Gr`�g�q����_�6t����gŃ�J��&��,my�4���m=��A�P�v���]�_+�6�IT��/;ϣmN����@"��[�Vd4�$5��R��r=��i�d@�%�`R5��g�r;��������LF��0��K��$L{��?�M��� �x��F��6 n0��!n��gJ.�"�T$΀�DM���O���� ��O�[�RF�!��:so"_}�������	�#ow���v~������_ƿa3j���WB)���!7����<��� ����cg)V�jO_u��x���i#��:XL=\�:���e�$o
F�1(���v +�ۃ�!�i������������Y�Q>(T��q���K�g���+��ý `������Q)m�ڛ����e����s��Y���ɭ��?Va���(�*��ƎՕ��/��"�L�D�I���ZE���x�Y�.�W��t�/��1�pH3 Y�S���Bw��H�A�yE�ȫ��z���<�lV�$9׆�stR���#����=�Q��=��.�B+R�O��O�g�;���؛�T�,ǽ�}�f<6��[6�:��,����U1��a֒*u:�@z	�Ң)�S�H��Wj��~N�L��z�,w����g���(� sG�UN[ӕ<������������m'�K^*��������������-$�����K�e�->2k��2��:��Z<{I�V'��q��@WwKj�m6�1���ޚS�w�rp�Fw��Ү�T�ɪ�>���zE)�=a�t�|{�Gd��eЮ��#G�+�
:T���K��6X k�3��5Q$d>���E��!T[ ��@ʓ�I�;�H�.�9e`M���WA�{�䨐w����T,sۂ.C5u�w�+8J+�v
Lˋ�s٠�)>m���V�����<��J� ���Y㈧�����.ag�y��f	9$�~+nD�G��7�x��`[�qf��O�k���fw:��GѲ��5B�d�����ֶ<��+�C�i��Q���bvt�U�Ƞd/�Z��v�V��7��O{�7�e���}l���'Û��� 3&�~<�Љ#Qd���4�~✲���k3��hNb��邉O�Œ�BD�ܘE���@g��?D�IkU'�-��#0���&eNB�F�=���%�;���E5���j�54��3Ӧ����ۄK}d@ec>�|���+�(;�C��r�0�����E>$0oh	��Ц�ᚚ@�:�o0��� R��z\)ɷ�$Os��N�Fݙg���M؏LĽ$d�@em,���Vh����E��U�����,?�h&�i�s�J8�N`���-��X�Ї��AI���ݻm�zk&�Ho�gQp
U3��T�)��E���ï���yНws��WaY���{vH��
z�)K�(#����1yv���4�TX47��O�ƚ1����9��e9]�S�!���b��������/�o�x��H�E�$��ʏ�e�~Sg_b<s��Wz^0+�w�O���u,�vb������w�f��k�{ i�(f��,1��E�Qw��ơA��鬡椧s��ZD�~̟h��a�l��f�c۳��f�+�����H�B,U�q{q�u:� ]��:��>vJ��-�=���	;�X� ��P'�U#Z�5����n�9�GR��Z�Q�t���`�ĳ;��I7'T�Zǝ/��=��:=�Fݓ��L�)��ݸ��y���,byR<>�K�<%>�@B�B�'� ���c�zou��.��j�o���?--��c���|����W�H�c�Fg JZ;�D�sO��J����HHzK3*e� �!T�3�܍�U�O,��I�d������߄ֻ8y.����h�e\������XI���>��wug_���Z'�� ��F�M'~4�`b���V��� ����|�������NO�D��[� �J�j����Sy�a�E`��9�eC���S��i_	yj�1̓ǰ�́'�Y�-�|:\�����|�A��a]� ��GD��w�s\A�f��1��BnhSN,I��ʽ�`���� �����п��`ιG��b�I�oo���F��T�/��G�С|��5���(�PD̕z��qu�2�����q�{G��)��W_��-Ã��˭)S��,Q& ��:�c� ��;@ｫ�<�Y��s�5�-Ն:�T���x���K��b�nǄh�M�T]/�_"�[��X$Egj$���B�bK2y$�O���=��_E~��NtX�U�������	l~�q�d��]~M)�z�~��������J��Jj*��U��>L	�3�ԋ��ރX�13w�x`�IxQ7:�k�{�^�6����J.o�����H>�&���Z�����EJ�}��}�l��$����-���@W�� "�[r�����	1��Zt��\�����!{�!���e3�-`���}F\B�Y,�,�>ןl�P�ПFؓ�zV�:{�q�t����Y7���b������/7q 4��������̛��Ͷ�>��/�G���m�A�3�iƈ�iLD�Pd��؋�@��{:}`@d�ݿM#�O��.�7�zY��F�}��[i|nc���vv]U�(��AE�n���|p$�#��A0%����9���|Q-�,>U��3��˔�=6КKx���[��x12!%���@D��:��C�U\�j�m��f�Q���NmD4�7�qjf[Xl���&�T�[�Xð�Q%n�z�>u�0�M�M�Gd�9�O~|&	9	ɓ�)$�i<Lku�Vh�|���R8J���:�LR�ѯ�Vr���<���)�4�[�rgS|����yM�S��A>�7�a�t�����L�6���������A���A���OI��Y��/�H6(B8�Txc����m�8���j�Ryb�/����1`�s��ţbJ�F�3��d���/(��򻻩��z|�~�8�R�qd�T�8�K�빿N����\j���3&E`��K��+�5{���c(�E�m�G��N����L9S���~���	��?�_T:64q�N�} �s����}\��	3&��xS������Q��<�� O9 H�t ���-�H-_�����EN�\ld�
���㝶�#`BwVyf�_O��r{ۖC�OAц_�S�ړg�Se^攆CR���n�
c� r��~!�"�9h넃B�Fk������d҂��%� �Q��D��Z!� 
]�B��s���[l[��r�nGe �y?D\�,K�Tn�L_}X#unx򜜛b��Z�SyO��)ݨm��H�Sb�������E�8�����l���~$1��W��^����O�^\6��hwTIܛ�C��A�D�i�D�D��`Z�TUa�؉��̖��?����H� ��v\F�A2Δ�S> �O@�NہZ	G7Kr�T�L�@��h����.��~�:�Ci,`���u�l骷�<j��cl�^�=VSɧg����!�����K$�Z�_Śe�>Q���D4��:8��c��H�_���e%_���	��Rf�v΀�Ќ�0����Ǳ�/��VlD�T垓A�Co� ���`3�|�T�#��oD�Kk��Bĩ�P*EA��O{�a2z���x=�C������g{���r Aޡ;�_G���M4��Q��kJ�J�K�2�@jϬ�Z.+���u���� �	u�[�s�8|�����_���Q_��m1&k*���7ť*1s]��w#��8�ǣ�JF5L���d>т筘<�X����Ȃ����s�t�iz4y��ݬL�ɒ���r�"цRv����\=�8)`�D�^�;��J��c	�q� *J�7�Ljk�G�>
�F١>o-��B�n�j�D���Ր�_�(h��gԹ
Q9��Q�����gʪ."�A't�kS�G褓�4�s=yeAɝd6��W��P�6����/5��F�TNV[��}����(�f�_d��)����>��
|���2r����|�ޑ5��:��q�H���DF�h��_y[��5.r����ً�9�MM���:�26�w�QBN�Ox�0:m��7C�*$���8ʉЊi��H�m�<jH��Wh6��5�4ͥ>�B���*1��y\Q1�Ǭ�����(���3��q \s �DP�4s	++|n��-ݓ�.iC���ez��i�__$o�5���f$Țy ϡ 	퓺�����A�x�WO+즧^�Zr-	��<Q^�NiYHP�=d�)!���4�xT}˖7n=W��ڙ�(oV}�P�h�k�-b,ީ�yz��e]�>'$�KwԞd ��Fۺ�����������e`r�T�pr�������D��W�[Jq{т*i<K3T�!��3�]b�G4W�5N5�5�Ow�9ڣѪM�nW Y�;b�s�c׿슀HmhrΣ�� �����E60�h����RE�l�˰���W7ȟh+�u���vdԜ�P���܅��Qw}s>X�fi��G_7\�l!�A���q�F!�׫Lm͵P���1+B�G3r+bF8Z��C5�zn�&�\�)ea�r�R�q�\w�\��k�O
Tݎ�|�@��4�bŦ��e��W�C�ա�O����^0����P��t����,fA2���{Y�l��t���@��4t8�2�L<nB��ZY֫�	}���rvH��ZFQ�[Z�Gh��o�cJ��f2�MT��#E�����w]|�<v�Q�8�ɵc���]�7�&2-�Z.c�� 1U^v���[v�2��.��7�4�l���$�FqØ=��|�2"���؉S��_�� ];��[��ޞ�q����u��f\��W�N�:i��̯�^�Q�}�P�2N�����R) .�ĝ�sԢh�h�U���"x��)lD7�f��|kZ]&��|=��?�/s���||ea<���Ƥ���C�����9	�Ex2짙3vKt�"���Fߗ3 �#��k5����*
C�����DϚVɫ�9U�>�x�����#��J�SJi�5�݅}<�~��M��

$��/��4�^]�����j�-�'�O��l���q�H=�����2��&e�ꬪ���'.�&do������#X�Ra��(�<=S:
��fo�_ ]���r�cx�A�]K(S���������ԧ''0�R�߬�'�I��8��YU7+����l��-�^*[�����xV����p)M7�F�<\| ��b��M�U`�Ϭm����X���T�:0�W
2j��?��_���C?�Uy��2Xt�8��@+~Q;D,(j���r����d�)X�h�6ߘ�X;�HHԄ�%���gJI�hw��abKʬݙu�����������RD�ຌ��&�a�[�f�k�oI�x�V�{��+Y������Hg���c9i]E7$�J�s�����A�]2�NFiu�c#t{���gm�v}4 �-�s-B#�� Tk�%�Aa0C܋v��bxY�=J	�m����"�����aB*e㓔�4ک�ݯz�
��[5�������#L�w�����9mWp�o�)�0�C{y],Ǝ>MQ�i�~c��711�޳���6>�����ԧdfow��	?d�9���";�#�ݠ��3F��PRG�F��)#Y���l�Q���*Ae��3���QXR��X�iJ�ɨ&Hj���:+1��m��F����i���@ ������S��䚆
tQ9gd���nJ���"�0�-E�ٵ\Gx�f���,�t��DD��<�%�:U/��_X3���h��JG"���)j��4�3H�6#�w����xB��Z���eҜ�dU���=4R=�U���9d~{�Qp�^޻z���"�c��3���w����o]���D�X�o���mW�K�R��.�KZF?kQtɭ�?+��-� ��_�I�)�bРN�r|I/i.^O��藤֖���~o���-���%ڻ�-g�	d��@�1�TLT������вν�ɐ�Nw*ό�	�iwr�|*�ԫ�܌��[����as��z�Ij]��`1��A�(�e���}A7D�5�����L��ٗ�+�tL���{���J�����%\F8�Rm3~�*�3`wB0�6�v��Bә�n���e�zN��]qm@��A���#��"�*���vQ$r�����z�x����@�K*�P �\�G}����6=�+;��a�lJ8���-��aq��D�R��?�:�%�0p~ hB��ˏ�}��ԏ�9���p4V�Z�Ƈ�D4) �$�yx���ߒ�,Q?��{ag����(O��&/0�k@z"��cu�[��߼���3���j��E5p�g�X൧��w�Q�y�.MC�g�5���xq�D���U3��@����PLѹ1k�^ 7֕Z%�o�#s���y���:��푉Ѯ#���y��:��S�d�7j��R�֖�|"|o�*^�W��˟��s����#Dk2�[�C�0���Dw��}�`'��[�����-�(���,H����~�0(�PļZ�RY���0V��'ӫ׏3F>R)���<�/�I���+a��"|��������ӗ�e�cD��A����]����xo���x�N��bJ!%� �d�)W��drGAQd�Qw��::�]k��8g�=��=����j'�&�[�Y�T��&��.�lm����9�$�c���T�8�E�����7g ,���҂3��1�?T܈Z«f��l��I�j;�$�|��f����H��]�\k��pq^�o(�:"��K|_^��B��ag6������y-be>O�=�ҽI|�����|��r�$�(~�ӾjK�^{�p��������Q8�ظg=,p���<���m|IY�[���ɪܶ��a�J@*�G�;�T)�?d׍��=&$bӻ�>b�����i��ʖ!�r���@2��S��n��t����32d�;ƀ9_�����Yr��"�6�j���yd֤�b�'e��#z�R�G�7���73���[��y��nlTl��a^-H(��-��%����RR�X�����|Ӈ< ��X�|���� ����v�@�F��o���o���H< kA������Λ,����;��4=-�E���t�WZ���*��,�Nc��]b� �V��swXwv�ؕ�e-(�6`Ʃ�>���ك5�Aq �v��2(�됟Zd|3���J�w,/iy�|�8}32�3e�߭���H��[��3���|Q;�`*���-0������t��*�A�7pď�S�sxq!�����&��l`&��'J��=�!s#��=������xK~6�|�胞����u��u�-Y�&y���v^��ڊV���w��k:2�bt����+$��IFgH��>���ї�;��M�ɟ�Shs� a������&V���0!U5�0�՞���܀��ö<�a�Tڕbs9E�s�l�(L=M8��ʎ��n�gǸ��M,wÅ]"��ƣwZqdsy�xG�!W�[��d��:�]�O�z<���-dD�.���O~�y	��!�ѓ[���K,<Kg�b��:�Z��N)@�+�ɐ=��ˁ����%�������7gdä��G���O�gRP褘�s|��J��/UMn����{�Ĳq�Z�}�c�9-x���K}��V�ش+��2�_l�[��.�xF=H�"�Z��~a�ѳES';ٵ��璍���/B�l�u@��{>�GAv��!&0�{��������y�aR�U��@�s]�7�'�="�49��ru��a�