��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k����W�z�N��V�?�ۿ�)t).��7G��ζ7��
�(_'�W ����T:�~Y�CZ0�i���sZ�`���Q��X������6x��Z ������Ë{Bfla���JLn�qI��s���sj���d)���p���4�EٗOK��u���F1ܱ���
vX�[>n;�&+a}�Ez&���"�S���}��Jm��_M�d���5�?�b�a��"`��׵X,���ah�T��s35r�|I�6�j���t9`�gӕ9XlҢ�CB� =u����k��0Q��~�0!yGHf�����_��6���������, .ʇ���l�H�Q�)X+��ծ(,I�������K�|R��!"�8��q��&�˘M��;�!��,��;���5�"?[*1YU�l͂����~F� Db�d!� �G�r
}��w[8b9Z��TTR�!Ɯѐ	�q���:�]���3��c[��et�;��N�w�R�Kw��;3T 4?-��,�Z9�r��"ȓ���=�9��`�C�G|`P˜�>�}�ݪy�*H}}���0׫�x�5D���e��b��ݻ��BDm0L�B��!�٫�3��m|x�Z�ҳ�=EQ[Ώ0���Z���tsx> 	����r�w�w���o&,8�>�*��K\a��t�~��wo���X�����zx�$�p$)Oi������etm9���Lњ����"����yi:�|�Y���>����i�+~���$�p���j?9�J	x[�����X-�<�;����αw��8�{OE	����̓IAM���X�4<�͸qs����H��N�V�Y|���#/ٴ����o縸ui�mi��=U ����t��M<�1�0L9�F���,^�/M��]��s�Xߪ��%h��)�t�\���D�Z��ށή�M�6ibǈ�����H�֣�n��ф�t�U P8~�8��Z�H�%<b�9E��4�pV*(��xY��d0��r�w��J�#;Ymu���X�cjr�DB���Wt@���X�?^�}75-M��� �ĉ���M�o��'˫��8��d*����X�?����"D�E�O�>��/�MJ́|1�ɶE$�Y���-
�������`�:;%����t`���v3k��&��l:	3��|��E-�(�+���I"���KT��Xf)B���rC/-ڎ._;��!hY{pL���Oh �,	����hC}M�}*�a����T&�6�bE�]1�R꠴`΅�t���<��P~"jd�u�r����g���WҦȱ$���aR8��p�$q��)
���Z�˽}nKY�7mô낛<P�~�cz"Fm�S@4ѐ"��P��lR�6�b�)�R�B3��(�~9px�w��=�o|��:%97De���xf^4Ϝ�e.]�J���7��T� ���댚nY˟���t+�����Hd��p���)ʰ��X��62�?b���7ׄGw�_R�����|������K�B����l6�	���z���a��m��3�)��q�\QD�v��l�����|�LAr�	�~�&��G�]�~��<nfH�)�50���+�Iy�*���Q�P��?���[r�?={m3�g��e\)��ם�h�V!���Gcxm�Si V���˙�& 0�J���Yzd�pu5Ey&f՚].u���X|�>&���by��量�+����Cﮂ�g�>�$H��o�9T�<
�H"�ڽ=��N[e���n�pTZׁ��ü��}��$So��ּ��Z,zmۤ�0@WsxP;`K$=�"J�$���^Ϗ+�xݕ�.�E3��`����"f 3��54i������*���UIgHd�چ8a[�%/�ʰ�$e��b��6�|[+	��D3�8�>�rB�}>�	
r�����sg+ĕ\�N�w���6ze��A��9�]baܧ��wnש�X�B�iu��o���>���%����O���FIzH�*޻��U�&`����ǭ-��o�����Y��.�L��{�:��;t#��{�5Z$�]�Qn�hw��@=�k�(R]=�D�0��h�ѹ^`���1�[�؇m��vUi����¹]e"��V&^�d:�?��M�W�5���W��B�$B ��=)�'�
�<�E�����[�e�	%��s%4�}�x.����a9'��˝�n0�P@�!7�&#�6�Jk��Mb�,�{{�B�L��.5͢�DK07