��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k����W�z�N��VXi^�p���d�����3X��#�����Hȑ��]�s��ތCdvc�2�k�[�E煶 ����#n#�5C�S�_� ����#'��pj�Y�pi�>�cZc��il��bf�F�x�\�~�Uj�
�<8�*�^��\���}�A$��I�?|/�J6�>�f���ƾ{����B�����j�k�J�3�"	i ��I�;,>#}��NG~j@7�o3>D0kvj�Z����Ű�+�>�̐��ş��E�iPy��*9P^c��Ԡ���"�ne��	�£k�)� �m毭ft�Ԉ�H��Ʒ+�i\)����6�he������H73Xq���Џ���o��x)�T<o�� ��D���e��z$��ޕ+�P)=;ڤ������%����r#��9�<v�b��4ή�9�nEG���W��փ�K��!��ʱ方2���.�]m�)���MG��h��6���h]�~�V���<�_�ǖ�W�?�n�p��B�.���¶W�u5���\܅�S6�V��J�((�)
��lh��|�xj���Pگ�Pp�q\?k[�xr��@���n���N�
�ʑ�~�UD�ο��;!�(��=\�;�@d:�� `�ğ��#c�����g���la��~:��[�H�6%�o>C�t�/4[ڦSl=�D���िp4�����
�����"_W�V�8GEn)%w[\52&J���;���p�]�W�F�H���lQ��:����ѕra��<�&����~��
`����ؼ=ג{�4Gz�Fǈ�b����OQ}�����<�t;���zT���S -@����,��d[*䦒p���q�&K��̞29��������j{��*`�z�x"K/�S�&��q�x�XcC�>��ʾn��"C�{+���"O�l��L�S'����8~��E�����i���D��DTT�sN����k�'�(������aqj:"7�	�v3/��a��.�t�Hｯ��齶���&���r����6��^`����^zM<��\ :�ݽ� ��K�HK���NϤ��jA`�I軟���]#:v��ڛ��t���PI����K�� K>��t�P�����c��C��(����c�-\�?�rJH֚Y��2��f$����'�їw԰q&���<���#Ͼl�h ���=��2l���٨�|�`��!+��F����̂{���N]!�	��¨<�q�{�<�%3�ݴǟ@��ϙ�*��8���hͷT.�Lk�<{9L����F����=��s��9u�u ��j��e;Y����;�Z#��5�&����ZB��Si��@��I�&k�DJ�Ϻ.( ��ndZZ�/<'�� A���K���5͘����`c���3��o��l��/�暲4��&s8�g�i��y3��;D�M酲E���uEX�#{$O�o8y�ucc2㪕O��d��I7�K?ԡ�6��@5VC�=�`Y�w@�r�Hy��h���~�. %�݋G�����P��r��p�Fx�an����n�0+י�	��Z��z�d�5�O�½�7Y�cC�"����ø8��(���d�������HB�*�N�]]("�#���� �
��eZ��S��;���I�B����v`Muz�7�蛜��J�,�:�󯏊<j;7��2��q@oM�,��ݛ��QR^=�2})�B�O�
�?N�i{��N��3
�2%�?r��sG�&ob��c��v{�*�x�"A:�x�2N�>�W�֎��[ªI�O��W!�d��K\r�P>�h:p\�������yK�v&'�����(��f��`/ej���E#�ſ2s�\A)���VO�I0%1H��W�����u�u�uRZC��uUe�z|�p���Z��	P.M���%���q�TQ��'�˙H�w���&����rY~����ܺ1��Co�
OB���U��)��<��`2IQ������|i}���_��vm�ɦ ��Ewή�;	I�:<�w=�@�׌
Q��`8YE[�����7����%�jO�t���/�.�ڵ�U:��:L��ӥ֛8L�a\����M�uD�0��}
'��q��t2]�B J���r�"�_9r+�l<�9v
S�T�*�Ǵ�W;��O�9��EÍ�	�\��Ё��c h<�����̡��f&�6��[�ND�K�}����FR�4��E��/d�5m8Hɝ��e��qۅ�;��5�M9���Z\�\�����ܐ0���1���m=&J�ss��p��lZmȿڍ�נ�0���9�b�M��)�@���܇uTR윲�4�j1�8���{�}@1p����R8M���<]��,�owt��5{��l��(���I�%�C?W��	���2�1��O���'r_����F�&��.��э�V��il����۸`���>;'�����'9˃�Q ��?t��%��.B���u��Q]k�Jڏp�:�ݦХ��r@�+����Mٜߪ�7)�QPb�D�ʰ'���w�Һ�gy�i����Z9j!z�2��>\)�#}���%@Āe�ƭ��m����ڳag�0�e�|�R<��b͔o}�����J�u�� /P���],«�q£ϝ�����������b�����b*���"��Uԯ <�u��-��^G!Κ1�?q��g��ؚ/��|��,-��~����}��T!���XL`��BCb�E�.�N�4��	|6J_� ^�����Q��Ou[]j��L^�-�y$�8K���ʜ��^�G�W�W��
?B�*y��B"�g<�4>U�Nٿ�pq�B�h&"1�{��FV?}u4�l�#�؍��	S=�5sQ����ȡ�9�R��5��Ѫ�J�Y9E���8i�Nw���i';�2�Xn��,�<uؖ�t��N�u|�J~2,Q�DP�-�'���O'����C���T�,�7�!Faεk@�L	�ۋ�}!Q � p�3�Z]���s�lX�,j0�(m��MWج�9�._,���y�r����ZV;*֣��Ө�S4��k8��Oj���Cp���d_)�m]�cЮ:��7��9��^�����'j*�.$�L'X#����i6����`��.ܣ�|@�� &�b)��?�&�oШ�W�c)����ن��<Z���e4T��wGB>�8��}�:�P��T`�����M�#�mI�آ{���cr�36g���r��z YTsa��f�yj�I��Y�y��;5Ŗ0���r�# ����}F>x��C�������Ν��j���֮`N�����j�/��0��������Xyo�g
w�"��wV���=�{{x��b6ۼV��R�=xlpq�+O���Dh{�B�{;��Qf�$5�Z�M��)�r�]$ݜ@�b	J�Z���᥺ف��؏.�Oe��ƒ���p�����;N�����
LU����ʛ�D̍��)�&�_��_w�I4\���!s���'5�BOV�sÚ������̎�Y\r�C���.�[��
�rԧ�YD�kq����!���ݵ�ٌx/��)�a\���`!}�/1E��:�-[oa.�*�ԭ��u����9/7�:G���d�-Z���!&`C��.4��:4;|�Y�E[���Aya��	,�����j�Y��J���^��̼N�]��և���)	��Վ�C���j���H}��ʐ%^Fu[TW[��w	e�<�ߖ����\�5v�O�����k���RkUٴ_�F�������"9,Ef\�Fa�B���Ս9��Mϩ�a�ʋ<8�N,V��$��Hf)���<��h���~A��t����	#th�i#�C�>�ڧ��O�v�ѯ�L�|F�ʵ�BS]�tÓ&{mZc�M����C�|��W�ҿ�;�m���q�9���(�#=�Ƕ�*�ׇ�b�P�*]ֱ	gr�.�?� �ǈd�v��K���(]a�+�ԑ���șL�ϖ$����i�I��-�!�B����y\�t��'Abm�h��TDI���X:���-�wTƁ�2_v�Sj�4�mmS�f�p�+�:�̽�4��Zc�[1�Թ�a�5*��O1B1�~�vX��}Z�ъ:Ɩ��J�rj'(��C��^կg�?"G�_7�+�t�����E&d�iv/�OӽD�Hņ����B�@^����O��R����Qv�T��d�������ua=]�.�~}��"!xލ��~���
ߟeB�h*�тܤtC$��D#a��������o*3�����rl�x��n��bK��
`^�ac�z#���/?���\+i���	������.��׍	{^sT;�Csp�Z�5c5�rkA��p^_�r"��f��^$�I��,�b�nO1�]��Y;���%P���qj�����n�M0�:��Wjy\��8-2QF�)�k
�o0/�Gۿ��^�����;k�w��oVS�K�L���8>ƺ3c)������M
��ڠ�k���´|��8�ѓ�A�X!.��|�d�F�bB�4�����ס����4Q�TP躨8�W���rщeL�Dv S0���}��G��1�}�]�����CV���h;� �*��ϙe��?.`�l2|���mN,2]�x�G9 �}�]X''
�V�&��п��r�Α���+�l���r�6��5��ƆU�d�z�]����aP@f�ݝ*�O'��)rW�Oe�!rEͮ�
��[� ��(���M�� ����,�[��~����)��5LyR����dZ��{li��[�k7j>�4yZ�*�p�!f�n�~zr�h�W����V�pJIb���H�1p�ci��x�	�ǯ�E�8m8�l��r��D�8�-jH�7>ɢ�(d���okD��I�I �4Z�F�}<I�4��e�L�M�J���_�`�Yt�Ɛ��#��iYa����E�R��uD�_ �_QV���f__����(��_3��w��֭թq�xB��)c |йW�������A�g�b��6_�b���%>�j7'�x�M&��y�����������0b=�˷D�'f�tn�������Z�-�.-Z�%u��y&RNn�VU�:���q��Qg2	�oZ؜�Z�?�������gH3���'I�5�03�k�;0X�YVC�-�M��;���cr�{������y$w�a�6��,���d�#M� ��Ș��M��!�f�]��7�,]��׋�6��:��L�J�ap�T�S����*jӠ�gԫ��<Ϳ�Ғ�x��h�@�i|AiuF_N����2�Ӷ��!��gbB�#w!)���뒲W�:A8;b8	������ta���Z�$�j7�.Nj�Z16A�'u����H�T�K\i�����sYj����#�+���M�	4ꓨ�"��Y�L`���z�بP1�sI������@}��������q�4��wz�WK�S�{ v�zS����_���a�ckDl�Cƛ~sGtN>؏�T����e�䉍��ဢ�	*Z��ס�C��Zd�3�#����ҝ���������}�x���
0��������R��᤹g�	:����%vr��ՕA�H\/��^�Z����C+6�N)�˝g߼PX���A�9N��c�H�0C��8R�9������.�!��<�ǵ���բD��v��	��	�j)���7��F��E|P�𩚇<��KR��xH���EF
�j���)���^@϶	�xѴR�����������?Wգʋ���%78v������ �LP3FG`(\���n(Z ���}\l��-Au�ֺ[d��-y�/�u�fR���"�FX^��1�~
��g�18ٍm+JI֣ :���>s��x����(��j�{���ǧN^��r"���\j�C����4}�j`��}���vV�tO%D��"�OY0汎
^{�����i���ȸ����s����4r��aEܶX֯�&��	u�T	D\e�F�o6���	G_���O���w~
�}�M��zg�h���loiW�P����zZP({�jڡ9�]��q�.����&;��PW5��>Ŕ�����inJ>f���y��}<�|6�P �
��~v�'�^�
�q_�����DJ��������`�ꖀ ����~zJ9���&"uN�T�wv������`�7�	�y]�]�I�ǌb@F=7A��/�3�
���p�<�Z̽�`�/�ʑ�9�G�2�����F�~���j;���K�	��e�r����)�����IST^����a�V��.�w<T��3��Ȁ!͙����ց�m��{]G!�Ed��6�;��?��p��A��p�����D�u'�.u:4gvh=��!�}������)���:�e���=��s�BLG�-e;��n�c@2�e�΂����
�I1s�f!�]��,ee-^G|�`�5֯og�? ��B$.������ng��v�1���x]9M��u�K6Px���L�/Bd,Q���]�
�hv�~�;�C�\L�;@��1�nfK#�y#�T�ݕ�d��S��I�>PX�j�+����4�H@��|��l�c,
���%�Ӧ���gv��ق+a���p�����b�m�W������ls#��^��$Q��������=,T���� ýfF�YdE�YT��v���8�7�fC ոY�{�n/��_� �VHPk?rm�y}x�a�U'~��Br�w��-�[ў�6G��wp*��4���+�a�d:hH۴tV�D�n������ ����.��F���v��u��q��8��D�O� ��
��Q����Wu������(sG�+~9��턷HL�A����Xm%�Վ4v/��.
�\4���✠T���$IAB����Ss'��k��_�Iv��x]ř[!�G�0J�Q|$��.��VI�h?�a{�H<թ"PϜ�8�7�1��9E8�W��r���ֶf�'�Dur! �L\I��W*Mz�5�I'�5�;޳��W�M�
�����=-�${�]?T������z2���_:����C��C���[�]f$9"VQ��f6� 4̓�@~OZ�۴Y�y�x!� ��t��By%'����គd5�H���cx;a˘A�Q�Xw���'�\ Ihi�x.�W��ST7z�m��j�1:˭��r���zP���4\�>b$�;�����Px�U`���*,li>�lֆT cV���\�Co��=����I����pnE�����)����ݛ�-�4�LJ��Z��Y�<���7�e��R�`_�K<�S2�Nj��o�������87������8���"�Lp�A��]ED��H8��M���*��J�f���څ��{O�k���+8l�֢�G8b���A{;���,�v���$0d��.˖PoF��7T�~bHT�L��nΫ��PnH&?1A�g��bĀ(�����:��G���Z����)���-�۔�D�6��U�î�h�NEw�Aj��E=/%(8;�(����c���g2��ߨX��Ĵ�ܖ���0��p�-l�'m+�HT�t	1'��/:_�'��t2�'��KA�	�5��Жp��W3s���Gtի��k��=��dvUa>A�����:/��j�/^;Iw:����p��DSfV1���s$�{Y�[\�O'���d��&�⎂�3��D�[\�M�ԬX��4@l���W!��ɕ���$�P΍F���b�w�����e f��=�w~��0n�(���O�r��W*� ]�e$.{��}�h�̲��Տ�h�S(�����ػ1��
���������؅o��,�%�lK�x��mcc�(#�9Rk�V�+G��h���v�R Hn
L�i=�����Y.�Pʼ�8�Z���'��{��Ƌ���+�q8�赍���[d�G̛�]祟,����bR~F�����݈��|����2"�'\K�HNM���ۇ�H��Ϳ��'R�I���?:�Qͫ���_R&2��P0�_� Dٙ�?W�.�$Ә�U�>��uMa�n���K7�;'�%�q͓�{|'�>��C�%<�/��w�������6���z�t�#Rf3�����f,�ԦLv�4���g�U�.$/	!oԉG���f3����nF�P��'&��j���k\�;?�kW`ןvr��ڎb�s���L>��%���=G�Z��b�l��<$��˥��'�H}C-��ru�}a�����P�F��(�ԁ?Q�|s��	b�����$�6�R�j�T�.�@=��L�f�3�nN�Sn�f +�1tA��ʇ{�}c�Xxţ}�\���=#̋�J��{#���`߀P8=2�m�Wj:�l����U��	���it�>?�%����^0� ~7�i����cA�qCw6#<�c'�|�
}i�iza�".}��d̤9�	�4S���T�/\�2�]��)R�e���j��~v�1��^�V�a�
ӏ=x�d�y�쁧��Lݑr�Υ2{��%��[��b�|�)�չ����l��v�����_O�l�zև�w�-���Hf��͸�(G=4N���s�jHkέ�ܧ�������@�o�g�ƪ��'?cj�Ԟ���W[�ۺ��WKo��En2��Z��F)�uY��&:.�%S��-I#��j��TqNO��X@�wjt�z��РGQ���S� ��|���~m�ai�S~��D���:�M1u�,@|�C6��]�U��C����B�p��ɘ��S�վm$n/�f��]ja?�[t m����*t�ݓ(�^>�T?γFQy V`R��L]�����9���4GE~ �nM$����J�E�	���,��O�U�R��<c��
�������_���)�+^�Ǎ�[�ݴ�⾍�2dvZ����;�KDGd,���q=�����C�L�W���KB�餒����A�&� i4�H��g�s�[�Mt{(�j k����Ba�R�)�ڢ��oW%ؐ�7�5��\��'*m>Y���B���As�l�_`��@��!��u���2���Dh�'��G�az.oYp���DP��^T�a
�t��B��������7;��~�~d%+@�Z����[1�?�cOw�����)nt��T�+`k~�~���}��N�x@�����}p!����^
����k.�5��hx���ؼ�r��d>
�!A��3.�W���5X�\����
��IZ��*$:�9�P���}P�����>��qQӌ�P�Ŵ��K��I��kdkw��&#�#�2��>�(����.*K���Yc�Ǿ�G�&,BۆEt1Y�Y�j��_���g���2�m��G⎶�2R|v��ʑ1�Ԏ�q�m<l����:�d�8鈥���<��1G���j\�4�?o|m^����{%��� 8V�T�,[����t�����nߙ[V}��n�x�U#D���F+��.��۴,����.h-&�8(�І����YBAg��6.xṗ3���!j��������͍�{��F>��r�(ZS��V���`O���F�I��T%�B�n[L�l�1�>_�؊�f��|&"ۜwn[�~dC���*,w�������zŰ�Tۢ���GYq���I�Iq�	�HSӓ'(����rU%�a#y�T�O"a�� |��iZ�/s�x��*<��"p{|U����������B�=
�C)�Yv�Q����MU�5�T��m
�L�>�̆�
k����(z�~/�Ԩ�x;\2��~�����R�I�E�VyVc;lс��M;_��u͡�B�E�2�*�4b��v�xCNCn$l��Bꤒ��Ҷ����[�!4_�ѯ���KTTRí�d]��v�*G����y�r�鳘�c ��`~��U��ke�e�c�խvk��"�%-��|?=,�e	͗T�����7՚+��TѺ_��\����P�a�M��r|��a8e�*����b�5ZK�.��B����4�g�k��A*���~�����;��!K�<���.��7�I`��|���o�ʡ�Y'�gkɨ�V^���Q���zg��/g���leml�jš�X�����r�{�Li�T9Ӯ���ӝc��ǄVdR�93�{�T�"5ߵ���؀����)r��,J�PN�-}�}��[��+��Z��F:�>����S����E:+ ��tu���޼���~ӡT�EmI��]4gu�?Tw�Z�Y��D�*�h����8�h��	ը+�G���
f�˯��xޓ)�ne
k��wI�ӡ$)�}�L�`�<������h'��Zx GM�%-��Z�;�Ʊ��ma�N*�4�!)$Q�08�z��Cu��J�T��}!>t�p?�ɝ`���p�/�&>D�$L��}�I\X�Vj��(�>�%�?�m���A�����������dZ�##���^���3&���i�����(�m�h��kx4U0Xސ7:7��J��1��a����_rj2�2mZ9�o|D��W�z��3�4 GX}2���=�&J��Lm�� 0��w�{B�S!v�N֨m�Wj�d��Ih.Z�A
^d1�_UfDc�!]ղ.�5��Qy5v,���r��v|��ҡ��1B�3i�P|�/<r14�pR�+%�$\{�n��E��kf��p�;���	bt?'���V� Zy�����B���9�?P��+I��Z/�= ��{�h��L�z�S��NI�*�yJ�`�³l�H�5龥4v�m8O�VM~TT�2�޾��,+.칊������Lԇ�̆P$bA�-v����Q���C�$�SO��@�^bw�.� 9/�d��t��:[��|�Hm=��\R�"�H��1fL��ٗ-f2��r���5*H�y,�,�L1z5 ��������'~�9yeYP��}�}N)fN:u�C��H*�
)0�A�8hL��\�>Q5��4N�˚�f8��p3)c�1�H��J�Aq�r���RvMޒ�囌R����r\�1_O����R=�$�3�t�H���	��0���:Q4W��}i�G
	W��M�]L�ʬ�	�q0^��j�$�H�`�?���]��sC��2��T̔�i���?PՄ���c��W�jJĹ�������{��&��
��.y{��?��M���c�6�i��9��>u���2��������3�,�`�}�~i�ڮOwNw}s�2�
�ź�s9l����_ľ�YG����*�)�bg8�_���27�n�k���}�Ge��h�o�s�k���x0d
`HXf�����8���ף��ll���Ɵ���eX���n�'�h�O-$C��tW.�V*�������6B(�Vl����ć+37�;�3��4'���$D�8G�[�G���2,�"e�@P�mDG��Sw�4���scԢ=��!��S� ��f8Ә7\�E��^��Y �g�Q��+�Z}���Y��CU����AW���'-I��p쿒�;�3ĵ��R�4���0��uű�c@E8j��dH3]�S>��O��	Z��fnA��AY+;q� vJ_�|�J��uͽ�m��Ŭ�P|c�t�[V<=�h��Gm�n�Yw���O30ri��Z�U�W�M��j�$֟z��K-a�y��uA-���A�
=�my�=�UHIZ������^�S[d������dDB��Fe��2��f۞+A�[��v�%ҽ�lLE�NOR�N�����ݙs��t:�p�b��T-���`�ҡ���Tµp�a��1�������%Oŧ���x�	�-{��;_�A���H���yG���s��[���QX�r���~�7w��_���ʸH~�̸�zF��F_c����ܬ����;�u��j����P5Jݖ�4w��P[��v�
:}�*���b��6��.{)�iR�t��t�f���wiq������N�6h#��m�����8��h�ǯbyB����c3�������+�a�U�e��1~"�	Y'�A�7-��v�/5>�������eϖgҴ������1��N ��ە�_��]��J�! ���~w�����ʨ��+?j�1Ҡ�a�cd3r�x�w�\�o�7k�9@��i���R�g����8x�H?=yM���]��H���K�ȥ/W�H�G3DI[��Ӊ����7��ĵ��:��A���w���X(��i���� �'���Q�*�J�Ӭ0=�t;�F�;eCU�Jw�=��c� �Ɣ3�٧%��k5�|�1�6��K�$�mC��/�B֒�]��_��I�i����!�_z5H�?�O �) �^hC̩4���5�G�R��C�칋�%�=�m#���\e�������x:\��s�,NV�|9צ���`�S�)A貅>�%u� 6�]H�\_nX����=���Dx�GI����h�ڹ	���˽��H�P_�}V��M��n����<� G!��㽅�J,k�n�G�׻��9b���t�uϛ�]5��c��by�`t%���xm匌��21>u��Ҙ_�<vT��P?PW��$E"|���yǆ�;q�8�	.�X2K�F��s�W�%W�ð�pM�"�a�ՙ7���c,�r��~�@�_s~��5�s�a�B���2� �O��;q6q���73j���J.P�&�=#v��I�r�s��?�p�q��+�m���#b�}\�E����������tUjό�4_Z�kn�m"͟�6�c���B<<l0_��h�2��<@'w�)�w�-L�d��I��U%�4^�$��Z�G�
 �p�G�9���N�D����	�t����Srt�ӡv�}^��=��Q Pߞ���1
?�K��#�(��[������@��!Y��*1���vTx�1���e��i��H�n��-�0��eB)��[��qԄ��)N0�^���gN.�d�2���� ��*��C���o�?�3i�M�����EՕ��z{���F�T�ؕ��i}�����(��7�}�r
[�u�����a�Wi�\ͷ��=��|��wx�Q��Oi��*��t���Ŝ/�XL�0h�����|p^G�u��y�N#x'�Mʏ7ޒ����Q`LƺB����/'�� 9��=#��hDT4*vcA�R)B���W�n�gA��"(��?J�����y���<�j�^���bW�C��q������ �����w�@Ux00�C�6��_��r�mÍP
���T�O��2��/lH���z�ãÈ�Ȇ^��+��,60�;OQ�V�!�{]�_N���a+�4��Zi}��uB�ۺ�^�F���T��x�'�����������+d�k$�ؤ0�.*���uEƺ�t@��Lh2��*���I�T�i���v�0�Ֆ�{�x�0��^��eVF��FG�%{1��|c<
��!���v�,k��b`�Z�K~��O��r�N����e�R�F2���uq��U�����-�>��M?V?*�������ٵ�\��ªt���K)9r&�ٞ3a����ǛO�9U����D�A�Nn(�H���������G��Z5�M�<��ʚ��c�ÿ�0�� �Ok���̮��z}z��T;YY��5����p�0���ʋV�q�����j��С��r�_�y�'n6�ΐ.X(dx��Գ=)�#�aP{�]v�{8(��(��=�v��g(I���ێ����E3�{����K��Yɪ�K�Ԗ�k�/��7@���13V�Q�h��Cדq���������.6��i(��;~ۜ�e7EUǸ<&BF4d���!�f>��å~�C��W���qk�ۉ���uq����,@�<6.��-*�6:�r
�ï�n􋒹m`�~ŁY���؈�q��B
�ָ��vi�1]%�Wu�*.S�$�C����kq�J�n����%��ڜ$���b��!�a�,[yw�,��0�4�vrMɪ�{h���a��
�3���c���e/!:.�+<#Ɣ�e���p����`�Ҹ�o�,K�>|ffO���zH�v I��/<Jn�A�^�*�ty$����������8��۵)�����ӫ(�u���Њ��K���$�cis���?���s�GX��o5<��ad�j	�:� w�����C�NN�G���QU)HѴ�u��\{G�?Wi�wJ����"��vE1��OŲ)�q�J���B�͛9�Џ��JJ|��� ���8�"�b��:mЯLF��.��X���^Q#4LOy;��m���~�IexÍZe@�q��Hp�v�f��\�;|����h�΂15���꽔�}�`쀗9J_MR~�Kf���-.�3Ǚ<����8����O��)[��'���b�E��v�"�`,Jb�z�����s'�|k$52�L�:���qV��Æ��@��QY�O9�;g���728�mxb}o�%���br��@QF5�́��U�w�b�h��۵Xl�*�ݠy�W����%)��ȶ��c�����pd��e���H1��q�!l����U�w���ٽ����%,
��p��s3�D���q�Ɉ�Q-((E�b��"��4��Ƌ �t�������:����OO�C���W��e�S��!���j�K���̭i9��"FT��P�x�uiRWl�l��@�L��
��r��|�>�ى�5"�o�O����T�@��`~�U�U��x�'�GT�*s�ZN�PC\2<`�C����>��Qs��̖�$��p�c�I��N��c�#��K-����d����=]"&��N�t1����x��[Nf�!4��z�^xS4y��7��= �Q`n�v��I`O!�P��8�& ���6А}����Wc~�Т�?J_iqͿ�N&c�]\�ʈ߰��/���s�̍7�$��<祗VKg�B��	e�ɩA��n"�!h�'k�+�lya��V����P�E� ����A�Rِ�Ԧ)Fe��0�1]��/_�JZy�r�6ڱ�Y�$S�b��R�q�b -EM��Z\D��G3��(0������لa�"9�������QO�;n$��gr�
]&���ZbKX�'�2h}~��'�O�*`�yI��7̽ɍSl�O.~P�u�%f�D�Pi֓�(�ñ�M}p(������%��%���**���">�3��B��v��%��_�dr�g����T�Mϟ[*q
� ��n}��º't�����,(���ɘ�@�Z��D�ZR�x��(t�莍��Y�ũin�v/���,rr;���	�f>�`�N�	���%M��r�vW2 �/Ȗ$���>mP=���waH��ۓ}H�xSpN�)\�]�5<,��4j�ׁ&��rc�,��g}:�W#��SM4�&'�:{;~
�J��w��g�7����,����j�g�:M�+� �����m�Ջ�kJGu0����aTc$�FK�9]E��B��9X s-�r^�m�_I�EU���|���/[�>N�Mq�kR��i����}��]�_�d��T�~)��qa��pH7jČӲ�F�s�_��.O}���m�~�I����W�G�m�C~O�l�4�J���� �3�����,���I���O6��c����y̲�S�#�B��+d�ˎ�;u6�
��gl!���[ӥ��f3ɇ44��5��M[o�_���4��f�c�F�M��H������7���{9UT�߄���c��fƇ={6��֎�s:�ڍ�e*�m@>�Pu 6�h4�( 	Qpp߇o�#��[�	��Iķ{W������S?�����V-JV��cg&O�L?yٝ�VC_�խK0�p����]�B
��$_�*Ք���y�"�Z��Hv8Ph/uMLZ{��!���#Z8fM]��um|h�$I�dQ: nt"���:^,�S;.LMfVh����+�L�W�B���ex����gM�������h~��|��~,���En�r��u�2�_q�O�����&^a��&�TϽ3le�Q���u���͙	~iKi�@	پ��x!!�f3���C���=0&��o :�dOL��a	� V��h\��z���8�&�&Z��%A�����ߏ�G�k-<̢��\�`�t�'��P��дI_?ˋ�9{�c���8Im>W�y.u�̓ϩ���cS��z���Y��c�T�4���L�nx��� �9�M6� bk�s�g�=�	t!ZV����vwrHa��k`i�	.=�e�c��zZ��x'�!m;��0
#�_��}��7��x�f�Z�>�bd꟞)E[����,[��)n5Ԟ,�0���jw%�,���[��1�� ��(��~�����o>'�,�%�
ŀo��7M�7��o��4{��;�Qg^5�2��q<�?^�q���?� [*�X�
�.LB�:g�7Ua��b
�S�l� �d�js.!Z�qHTXj%����pacg�*���Χ:�7{;���m��#��T%�?�Y�Mm[��ַ�[C��*�!�<ҩPag:�Ԏ�;�ǻ��q�xRX��2z�����l��^�A��p]��/����+�7����Oro2�B/�� ꉥ�n�:e�H��n}3�u:�j�S�!_'e`R?���X�?�,�B�4d��6C�$�)]D�/�;�d7xV��$�[�l�FԴ�p��hp3�ƙ9���^����,���PXZ�Һ�-�E�UKN�l���v�+���ͬ�ݰ���|!�t�fo��zt��x��CL1�m��| �i�ve(|ｦ�f��(1�D�v��VVx���N�h+�c�%��5'+�Rf��f%�Wz'��f p~9�p�W�1=�d(�	h���lD꣚�a�WoM*�����ys���@L˿5�t���\S9�8����u��)��p�#�&�Of0���wA]Lv�ƥ3�ٵL�Po.�M�z�S�+T��*��;�h�Q���a,	�{��:d/:.6�`��z�U��3��,L�Ǻ7N�9vG�	��E$֬��M��(f�=�b*���1(��f��^s*b���!�Ȣ �{nĴ[��;T��3��3D���e�=q��E�<Sf=�sbHYჵ�R��4L��)��Qe��C�?kf�
dZ�,�2�����T~eNm�L��g�=��H��.�r8��0���{P�8����R�tt�b/����zr'�o��z������������w��v9�ϑR	60g!��)Q��(E*�0�V$M�WL�	"|1�-hS��U��f3�0S���@����$�2Du�0�YYxkkC����n^(�3�U��u���A�j�AAA��-�I�v�]�'�}��i�s��	��ą�Guk5��]4����� ��j���h����F~�l�Am5�4%���\����"f�׸v_��a�Fa������ Ο@��_P_y��2.��N�`Xg%�@�%���* �5D
)�z6�����4�!�F˳��9cw�牖�8����I��g��o	$9�&ju�Z��a܈��� �尦|�۬s������f]�6(>X�ӝ�����t�����޲�nI�H�`C��3�p\���t˹������\�wm���nrW��ҥ>J��{ �m,��2CD:!ؘ�
��v�������d�|ݜޛ�<�u��'�&=��^N^p�N���c��r�Z�e�"c�H`2m[��y9}u|�;�����i�t������s(���?<�G5�;�h��V�2�I�7��7����jqҢ�ɝ)��.����ǭ�����M�Ǟ�B5���_��X�h��Y��MM����^yd��!tDېϰ6s7R(�������ܝ_�}�$Y{��(XjiF��]��yH�A�	�	U�T��˫���X��˪:-B��;9�ݽ�`z]��H*kpc�/ AO7Z�p�����)��j"�e�u��?ڍ�ܲd���u���]�t:� +��kdA�-ń��i�o6"뒪��Ö5�
�s���� �:zw���SԶ	`��՜�e��>�U�S˖�*�o�hs'�i�ȣb(�ix� o��&e%_ ��x.XG�P�#��n�P~g�T.h|z�NC%Z`.�HPgL��a�)�)c i��^D6�	0_$��+�X%�ܑg��s�Z9�X��E+��ͣ/�hݸr�A��x�0͔�)��H������MtO�O�R:à��ɱʤ�A^7	�wC!G�2�����JVs�E�>I�m�yb�_����Y�.D�4e��M.�1��G�C��ݛ�e$N�p:���u&������1(�CBA#��)d�%��oT0yr�7�|A��Y��ʍ�B��(��Hg���d�t[���,�1g�,�]�q�"�뿯�K(r9ׂ&� �<�
���� e���l�9|�,���<��7�Q�K�,1nf���ۥ�/�"g���LO$�޲5Ҏ�9'�9���/7���E����}��G�<��BM�a ���_�Esh �sQ)�1:ǿ.�,�S�Sp)��d��7�ab=W�ż@��4-���@�>��Pװ���Ľx6щ~&Z�FƓ�$���7g�aeO������j�:��D��"G����⠁��%*07N����gQ���m��~��J���S ��"�����X-�$�D�9uw�ѐ��U�}�k�����᯷p�rFV�?8-���,�E7O���#����:
z������r��nt��$��� ��޹+(�h?a������%䨯���Q�oL�_�K%���� �J�u+��<�F �.Kg�!:,�"ian\˓����пȕ�hk��G�C#W*��x�~n)SRh8h�!��HyĴCMe��x%X\4�X�&��hw��M���.��C-=�h�F�н�l���ͷ/���I����.���I:��b�&y�:g��	8�!c�ߏ��\ T��A�Ŏ�U�Z��������������s��#�^,�Y|znc�qݧ�7>pH����"��>��f��_�
q�)��r�x�+���W���
��B���L)�?��ϴ�N	�⸸�\u��+���=����AO��x����Pۻrf FY��%c5Cli�Dv���yP,@:L^��8%�73�4G,Du�W�zʮ?��*$�)�?�%�	��.��f]*��	�(�m�V���J��]��g��Z�]�����}%J�������}mr��y·�<���L~��?w��� KtS���hA|�\�SƢ�ɦ{1�+�͓n�@)��k����U-
Y���N�ʀ�lv��hB>�(�U+(�)jC�w]��Y>e��T��!�Xݒ�� �tM<Cl- 5�5:Hp-^�kAl�3���?�ai��3&�"S8NN�-$���[2�������^���	�g�n����h���A�[�ZN�(��D^�i���4��͂_��&��ˇn_�YYT#�����E�7�-1B)�V�wH|�V��j���;jc����1�SXp���IE��[�~��q�F�h�f��'�Dr��+�-��gG.�9��`��t�MI�~�ÿ�Ds��}C@z)u6ӄ�Ok������wP#s-��D�˺z����n���>r�w�O�t����:*�_�l��ۍZGؿ�ȥ�B)u:t2JC��
����{�+�;s��{"�H���=ZclM�Kur�f�'��@�)vx)�]�/�	�m�l)��ާ�����:	�� �l����9��z���Z�O�V
�< �>|����"�]ǈ���&� �ȿ�(&pVKhR������A�D[�Ʒ�}��Ug�MT8Q�e��c����֐G�p�X�$�3X��.�E��C��[eh���"F}8��^J���M������:���'�Q}� Q��؄Q�1�7���oX���9�ʄ��̐
?�e�7��r�DG�\	o�W�*�Qw��5ys{s����(��+M>y�x���&�y�t�(;��F�̩i��T/�Q�yfV�\ �P�5�E��6(�M�u[�1�s����O�M�����/J2Ԓ�m.�(��%:�9H�!��s��Ed��xL�Lr!����F���Q���%����GT���������dn"=k���p����mՙc��+"�;)��Yd� ���ќ�j)!u�~�%�ט�UI���qV�:ե:�dU����춌�BcC�4��5Ƕư�Bزi(�N��gIA�+�-؆ZC%ޔ�ZD!�c���_!�E�N����	n肂,T��aq&ͱ}���%B)W?x�����0$׈�l͐��Z�8T�^�����z7�.�֮��v��Q�y���	�(�4�l����J�d�1W!J`�#�E�=�k/��,Nqn��h�(mp90��V׆ɏ-(���gg�<S����ŘadOmx�Qy>������Tʠ4`v�{�!p��;B���b��)�!�,&�]�$���X�3M�w�	�gH����ʤz
���$�:�(�-D��g ��r������Zk��k����{.�Q�C��FL��Mo�?/Ҫ8,�q�&q��9��pv�)�}�|�ӹ��Zazsʑ�cr���3ecV|�@ 5�.L��q���ć�T,�4�m��h��%�����;�;b ~HI�W���n�,2�D��"����ޭ��0�0:��7������7n�>i�dv������t���5��	Q��HDA����B�����!�J )c)�e%AT�
�H$Q��5�>��Zש�Q�CX����<���M����f�E	��G�K�i=g��%P����=H��	3h ���)��]�Ц�ȡ��!���<����֪_a�qu���տ�8�n2��pQ8����Xh�1�����d#p�.'3`�%Dl���Q�<~�E/Gv�3�S�`Y3��S�倒��(� 8�S6��������]��趞d��an�U��\���$$Ѯ-��c�Χ�%���C8�r�&���|a��սM�{�tJ��B����3B����m7��[ʝ����	`G���z�2=xEk�6."�(-�m"�5)ɺ�b�����0��^�'\�m��Jq�n�bb;���'�p�'G�����?�����\���̯�s	i��OO�����4�T� �l����5Z
j�A��!�n��+u2"�#�%+�$�A���G6���-���	ˀ��8`����SN���7�Ҝ���o�p� ��k5x�~��9/��a�w�������A��LEעv�q�1p���� �ݍ8iK{|2�r�~��c�;��=n��;�4!I�  ����ۚ���Īd�k�J����N3,n�I��X��P���`N�w��ڑM�u�q"�v-̴�d5�v���N�K�D$7@����]LK�ڬc0sa�~�UBPa���҉D#9����e���C8%�S��,c�'_{��?�H�ƶ�b���!��	�vI=�}cD�K�1�T(2bi��Е%l���=Q�D���zx��AyG��� Ŧe��p3#(1O�Ml�#"��i�"v��AS�M����-���t���!H7+�Mƪ�2��ġah�$s����A �0	�a��ҁ�͝���(\�@&��#���YȒV���L
+��D�rEl>c���]�P�͒�7Hz!��Lw樑��I��yQ�G�B��j��I*�YU�㠮�f��.��5�3��ߙ�g�tT zO�Y*CW��%�R��_���ܶ�['�r�C��'>�V�c����N0�8�Fg��%���y���>>M����I�@MatB:��dgE�jC��,��<)\Sn��t�@Hd���.D��m,��b�� �/jt��Yth����Bn�-��z0��4��s�����(� f�2�fF�EQH�^���=Н�&�r1��Ɗ^򴱬�7�~[b�B�P�|K���=��7Z�g?���2>th�'��@U&��;���S�C��S��R���U[��C?��R�Yo�m ^�;���H�ʗ�5�=5z��8Waˁ�[�VI����E~�pFC\`j�7Ẻ��&[��h���2�������rP~�Ԙ3���e�����/�W��,�cB��Ix�pQ�H�	�<���aN1-�(���]��ߝ�6f}y�zuΝ�{�HFŰ�H�D>?��D%�B= À�>�{���CO������/��)�4.�Pwt�W���=�8v �)!����
؅�9.���wO����X���	7�Ã�#.Vpg�Q/�z�~2��fQ��=l�?Z�A����;�s��o}�Y��B�#�!�vcbh�O�~,?�|�[Pn ������/Zaa,���b�GK�\�U�M����NK�<f��A5+�$���jZ�3����F$uv��j�VO$he' �t�o�P�E��9�9������o�Z�����(��(U"��Pi�Z۩؈ue�Ǯ�b>�F"�(�o�+����C6��T����z���=ҫy���$t��g�^�Ncn��@�mx�҃a�'�,�kњ�?fˣ:��EH��zj���u�":Ħ){ρ�U�G}�:�DW�Pr��y����j;�RK����j�a���b�Û��v��ĸF	_.ä�tc����Y�5k�1d[�1%��4��>`C�9/8���M���:\-����΄�=�����f��դ��A�<� G�\��G�1�*/)w������̫�a�E�G��(Ɔ��1<���W�-�i?�xU$K��3D��<�G�L��ix~�cr�,�;$�r��,��}�9F΅���mFռ��kF�0BV|[��[�_��U�k��K~&�xѮ�"���ztB�vW�)7e�1z�\+�G�n��Ћ����$HB��O�\���M��s2�0K�27�Y�J|D�	�u�x���7�� �̦�8l7F���)�#S�Ȧ�F���\������b�I����9����$�M��!;��7r]��:�_��/#Z���ʬUY���Bm�Ԙ���e����gNP�<�`s*�Ubì�1d^�ς6	O�z�p$D>ӟ�#�ס:Ӟ�dΉ�҅�#��J�)�]w�E�yՊ�̤rt����譣��g)�U�����!	؝W�=^�X��xUN�#����m�E�%/�3���60� ��2v�aZA��f�����@�U'�Xt%���1L�Bn��ruN�(9��ڬ}���O���Ҷ�����9�Fs`�gяvdS�A�7\y����ȑ0p�ĕ�����Ku��t�6'���:L�Q����~�>�#w�`��Ȝ��y����/j����a7uJ�|�]�{��i��y�'�ⱶp����%p��8�G,Xr��v74�UҷU$6w�Ո� ��7m�V�r|2b�&@��m��t�*)�6x^K� <��q(�픗{9Z���y�:�Q	��L�>{؂ �h�Y��k�5�-'��4"砽��g�&�P�a�����o�i�%�����'�T���`�W�}r� �w�`����|�g��g(e��>�p�Yg����F`w�QE��0���y�Ex�7[�u��qa�P]M3������v���ɧ5�0 ��7�3���C!G��(��<y����|��v=���W��0����v��@����X�~?盱vI��[ d��Z_*�>J�#!:�9��ގ��?�Bġ���͠1�^�.�
����^�Z����<t_��Q�D�C� {3p�nO�ͨ������u��>O�w��bt\���ҩ��#�x�i9�	 �˒I�h'�;J
��4�)�-��H݀�ٷ��D��p�9���q:(��7��E�(�����n�[��()3fx�᾽l�T��p���Ěݤ��C�s���Е�;�������!Уê(�T��h��ν�zU�����0�����Ƅ���P�ҽ�)މ�s*��s��r����"��=���dK/)dR�Pba�g�*�L�F+�*�3Z�ԁEg��p�9����%A�ֶ������h����͒��<߸Vx�K4I�fY���>&lxOX���D���0��S;?�Q�����2]�i�K��$�q�.f���!5Q�s��F����/;��z��������7����(�]��v�xs�3�lk����8�.�uf�?ߌe'��-	���,5V"	S�/,�F�ue��3�%f���Q����z�' ��"ѡ���G�=X~��i��}�yV}U������^�q�7��>�Zn�#d��骥Z|���B�G�-����,ݵ ��q�>����v�#�6w�[��nB��.� �MB��I`����?��#?���rMf2�XǹC�Hhy�cQ/J:����m�}��/�� ���-��1魎���c�.9}C�ϯ���D��Y���@�~0Q:������"��Hb-I>��P����1Ǹ��e�5 �~�
h����,�4F�^l϶�lݨ.ƿ��ӥ�Bdt�����?F�b�xw�Rl�L�-�n��+����%%�����/O �Y4����F�	��L��C0�b�,��qh�@=�7���{�R����&�ۻ_��lY	I�g_���J���|
��腡l�c�ʬԬ�<鷽���v��Y��	(O:�F~	@��j����<xz~�1BpeM`�M��0>�x��ttZ���'�"����=ց�������D`��V��UO��H�=Ң�����c��	�;��gؗ�d	l=i��9~�LWh�氱�A�\7��*�&F��n]��>�܈�$,>�9�^ş�����:{����]B����kJ��H��w�����v��0R�C�p=��x�X-<1��Sz��:��	�����m����6f����-�e��u����/a%�	37,��m7EI���$�n����tAD��ujT](\���8�E�كD��Q%��b�x��N�ːnK�n8�빉0��m[ �c�L�y ����Z��������^1� ���YR�X���A�?{=�.y~{���f���N0�n�:��,,~YQj��6�\�?m��E=8�M�<�xI����';��R�l5�L��P��j�$u3K���V)�e��3d�����?��ǎ�-�Ӗ�H��{#'��q��ċ������I\��:έG���O�4��H�K�+�;�L���Yϥ\���D���y�R�Y���۲�=0�be�$*8�e�%?)\sB�W�#7��!˱rf,NܒA��\�c��z�E���Ƹ8bb(O�����$�<�	��1�-+���c���_���KL��(2�+��:�I1ܲ͜�N����Qe���sjk8��|��J(<�(�++~����8��*�)I&�@L�WbUl��e֜�S���W��<A=R�ե�6_1bV8b�3+J0*�q2��F��[��c� �%>�7��wZ�q������D ���O!9D3�~�ő����%���g J��z���S���� �ch��{�;�pxEH����f��sf��EW�s���o��Q��Pg�a�γE���`u�'��"B#���N#%���,6�ɉ�Cc����^N�	N���/Z�
��5ģ��< ���Gr� ,%��s�����c����y"7*������S��N�����dh�N��"��g@(g	j���f��t���ђ$�F�O����Tȴ�
��Y�|��uiӍ��NHzw-X��>�}\�z̰��K�e��s��ȉG��Q!�}ƭn�+��W�y�m���ig��7��������l_������#���y��s�rq;i�zx��E_�{К䁷s�͎1��+;p�k��8J������{m���h���!�u�����&�ꄮ*�A���
��:t��[��X<�Ls��;*��?��nf���ք&�S��t`��c��H���[�)�H8�c����؈�E�����lu1��PY!7�L@"yw`B-f�kQ"j#�jHm���!�<W���h.LN���G�fU�y�pg�x}P�Z��0��>��e�����7�Bc;	1ܜ�mwA����__�P�lB�\���,=��	Q�����\v���2��0�C�|�2�)�
�7.�؞ܛW`@�=6��Ao���<ƨ��#�t)��Yq�	�׬g�_b/Z����yaV(Ժ����5s�N�sB|c��V�x��%T/
%�dg�$DUac�/�}䟠H�g���1-keވ�~Eʖ!�?��[��_��Iaӎ�I�TB�߬�Xm�U���Ej��~�]<��!,\�d���n�' 
�~A�=���Ά,Y�\���u���H�������Y5\�f#R%[2B!���!J�/N������$2F��
ㆫuO0	�E>K�5��i}����,�'|�N/�<������n'4���
���js{U��
�ss����i�$��.�o,}Q����ff��#�