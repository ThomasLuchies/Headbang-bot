��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+�������;���ȹ�v{2� ۝ߎ#�W�ӂ����ݠ��>_g5���t͉□K2���Ec�ſ��`\_��cW��Y���NB��*�!�#-/�����0�����e	�.ZDG����g/G�lз������s�VS�]��	�_,��ܳЅ2꩙Ō��M=룯+�&HfUk�@��%��.���cm���pZ�^�&]C��l�QQ���UicM���*�qz��ZU�^u]�2�=>���J��מ�#�^Ķ���l�\*l^���F��A��N�QI�������T�xĞ��pǚ z���4��)�7�z�wcl9du�f,u���� OK���ي�H�I� ��l��.O � F�		�,& �����ͽ�`� 7�(������,\��S�!�4��ݮW���l@����1`q�f�>�U�g��E�����a�md������N���+���+���}���t�
I��-�&���I;c�C&�Q�J���5땕�?�Z|D�YP��e�|*���#܉B,��S�(����L���͙�p�&d�d�d;B�Hᨷ�ǻ��qa�+���  YEɃ��)=��������Hr߈�/G�S�>������`0&	�wu^+�#C)H�C��f�k��U�lv��v��״KOgC�Ѯx��X���8�xh��]�
�J\:�68i���Z�O	G���[s�B:�E�6M�x=	��Y�hw�946�֊0�緪&�td����q��)6�wqx��L53e�ș@h)�}Z
{�z;�L� �HW�o��>�������T��Ք�x���W��#�϶�s��B�t~��%B8��S�96C�/T��C<����!���:o��T�v�3R0`j�>��V阜��[���EU��J����dL/t��k,`��:RJ�B�I���'�9)�@j3VӘ��Jzxf���:��t�	��-(ȡ(�7��96C��Y�S؝�&S���uK�	��z�S��U/* �1����n+�����2�'����N�s��,�
���՘�|�C|��ۢ4�"O[WO�[&
�|!8��E��y�����#	h��3(�YZŁ)�<���T�^R�<�{�PI�D��Bs󎋰��mn�=CSw��I��%��������21���T���1$�n�Q)���*���i�0m���C
�dԬ�'���T��o�@���@��n�\}����؂��ǳOpΗ�A��q]�#V&��)5��e}'d��ʾ:�?C
��[]�H	�v�^F��2��V��+:�K�Q�q4b\����I�������D; e�H� s<a4KC�̐�yAÖ����w_{^-ԟ�+V��s"��*
������~37U	���D hM��%s)�U�����K��-4�k2�ǧ�k�C�t�KKři�uI�M��.0Yc��eࣶ5�*�e �DmU�ͳ*�1ݏbun���n�͜a��@��i{#�(�w�{$�C��]�c�t���zGY�'ά��fv�F$
�ai�iv<h��W�Kh��~�6�>[�� �q���R=��F�c��X�p7��ߌ��c�>X-ff{�u�/7�������b��{2h8��[F
:�*�>)��CT������A�K[�i��XH@�i�ƕ|�Ǟu�D䝫E���k �D�U/�2�U��Z(vJ� �٫�T�&xA�����!U:�5,;��;Y��ʓ�<2ϼ�$޿��\�]
�w��^��d�b�άP�χ"�D�r���x<ŧ�>dbb�ʐ|�&�8��2�4�Or��횃%9����2�gڲ�~�V��t0�V9�Y+рa0�ʣ�8pk�^�Ag������Yu�@g$���P�Ѧ�R��@�U.��Pw��a��IG{�c��:m��hW�?���c������?�*fP���?+��F�nN#F�%�Rd#��Pi�;;��6\���[�L{ b�2�������BHj� _t��V;R��z��@��*�٦�1��hR1���7�UԠI:�7�}�5�$�mX�aֿ�K+ ,0\�b_h�3⷇0���v�U���-�GH�h*�.����J6���=+�d.\VtXY�Z�l�����iE{PܤQ���;�e���"�S|�|2�F"�>���3�z��0���o�vY��1Ins_�zF�3�~�x��JPX��?�(3�7���Ik6��[m�?P5�.cUQ����k(�����mEE=���K�9L�����C���Wϻ�o�c��X��G�g��A��lԮWk�F��YjΒ��w�>����L�+\���|���y�'?��7��.;Hng�7��=��D�Ŧ��gn��iڇ,1A���}V�è���ŧ��io��u�MV��bp����t�AT�	$�������� ������u��Gږ�+�X^a`I���9��/�O���gy�ݤ��A����YG%��5$��璵�b���/�bm�^���9_�����{;�H���u����[����Tx�O꾮��e
6���m��3�m<�%z	��߭���ϱ��T̑
e�����~�g��Y#uo��myG����Ϧ��|�ِko�X&�Հ�;~RO�n̽�$<R}Rv,Ou��s�ذ�V��,��������-p �f��`�,��q��~��ӉX��x�^�Q������3`��Wj.�>��=�8p�4���	����N�ڈ-����y���(g��hX�|�P8~���U����q{���� ��7V���9WN�Hp �q���R�3�!ܣ�����6A~�S�dKϞ��Ы"�E�:J�����B�E�����zE^�V�G��mLVH�R�����It�(KTb��� x5؊j��t���8�2�ױ�H���EY��Zl)�_�4�W������1 �1.��خ��N$�wT���EiC�A��
�0��t�'@ρ��ml1��s�5��	�ЂJI,M���1$�|�v�>?N%r�Я���IA8˒�3��2���_r>2��$���0w��݄6���[�|��o���1Ϩ*�x��P���m��k6G.�0�o���i��,���Z���{�wK��u���K2�5�:�)홦 +%���l;��:a���:���b8��}s�(�'�Dʻ�ss_}W�^]�0���F����ϭI�e��ڤĥJYZ�Z*��w2��-�r:)[�J6:���hi���QbQ�Hs��*�v�
 UT��	k,y3Y�tn_u�t���`��q�3 �KHk3!�n��ז������Kd6��xE��;�V0,<��X�_'nh���|�����1Y��e�?G':��OY����d~'5�b��<Ww	;�̫G���
d O��dHȪ7�Y����Mf��g��r��e��@×D8/!Y��n����'�����ŉ� b�Žt!\mwl�����]=C4���݊��̀��IVI}�����`�6N>^���x�M� �?�5��r����g9��u�_%�@��i��m�p�;��X���0z���)�{��]�O��X���\T�T�Чm*��@Ǐ�8׾s�w�<�;z�c���J�='4x%�Y]1\�Ʊ0����|��6�P\Qfَ��Ө��.g˳��/4Ŏ��²�V�)-��c��՜���\M�3V2e��}�P[���e�d{�%1x�Q���MQd<x �Hѧ�&N��\��8]��e>��M�\�#�2����8Й䣁f�E�4�:���Y�����I�Q������v<yJ/{�-c4�iD̐j��� LN��lql@�d_��^1\��ͦo��w�P��B8�����x���rnJ(� ��9�M�J	��A�1<1n����y�K@�am�P�_���Hx��B�?BJ�ޚ�%q.�tBW��/K\gYWr���T<A\�K����Xw�?�p�<�{Ds���3�!��f�f�<��y̱�i	�칼>i:#��ݫ!��B��荩<K�9%_x��em���H�Sio���fIO�.�O��5׶�wVZK �$�UR
Y���$�2��C��`��z	��7�j����a���Mz{�����NmS#�	)�����DiZ���خO#��n���������/��
I��H�Nl��E<�RXG?l����Iv!�Hj�e�k<�K)'�k��ҚX�	��>�$7���e*������7���(��S~�����~(5�b�6Ò&2U���� �s������.�jF�j��] }#��N���T��z�­��[��`��3��`� ȭ���Z�u(謷IqmO�:$���ͦ)W�O#r�䉕�p׺�6���qoZ���,f{& kS�\C�	f��D~�ݢ����.����8�df#�.�+kF��°T�0�9�+�/��7�!'�ؑ�ހ���d�"���p��u�_�`�{f7a�
`~����W70���M|C��7:^9�����ƌFۇ�t��C�xa��o�pkWV%P/jW�_,��Z�[%/��AM�@�"�{�I���t_KBk��u����]U�Q��&;���fބ��u�b��U�~h�yh餡�l�CR�!	t��~�M����U�"��-�z4a:�Cz^��WAL��s���A��	9�M��)\��W�o�*��7
�
�`D{�N5:�J�[��?U�^��1�h����MʴǮx����.�hH:��~QR*�Yw� �T�w�41\7�+']ٍ"`Xy�%�Z0t�J��y�R6�?s�q7`�&?�ioA� �44�)�c�m�:ϕ���^��<&+<J��[ ��p!�b��������\�y�r����xa��6�ژz�à�<K
_xq�e'�-Z��
G����/3�:8�����ԗ�Uy�<�qQ����*�%6�gI݅��d��y���_�;\ ��Ҁ�Z��mW���{)`�U��A�+J/9 MGs|f�4��l���
ina�qF�)��U�R��hW>ʹ2n�)�R�b��ղ�[��T7d
���6��K�Qiվ�&�WIQ	������i�Q`�Ww�-*V���*"[:w���FU���@tB��S��������qR�w�}y��\��kɼg^�L��PP��&�Y��!1����>��9�t�d�|G���1,ɊS�B�^��|��t��F4����{U�J����2imk����KHX���EHč��o���>�ٌE�	F_@�~�.�p��:=�*���Y/����_gf���+}�90BCҲE��"�#��n�=A�s���r�Y]��#v\�8t���G��qD�[��*����kp��N�z�׆������p�������أR,���e����{�]�\����d�Һ����� "hk�1d�W�� Hg�͓�"X��`��t���R��&힉_��y�:켛�����sA������e���8����p_�+�a��=���v]�z�/�b�����&�v�P~�A��9��=|����u3ب�S�����㔞�^-�a�rx���,�.Y����.0"!*դ2.�h.nw�i�~�?�Ϩ�%��fM�Y�2o.�����1sĒ�w�x�e2N3�1^y�R6'Xշ:����fo�	��.�дa����B?�o�{Xl�S�\e��b��K�6�p%cϻlq�*	��,�^K���B8����0��C1��HV���Vٗ$Li^�DZ�=�V�3 {�o[b�e�M+X�#�4MfUtyX�������^����{j��oQ�Z�����c����-<�����k��1�� ��r'1F���ѯ�%Ԫ�'�Z�3v�=��N� ��Lp���{�j�e۞������(�$��)�fW��8���X$&�\š[X�S���S�	��³D@y���4�u&F���]�}v�	bjR>�Hv0��e� �x��U�9����OKQ"���鹦�~�,~�(2f����_���4l�oe*�c��o9��jh���f�Ko���Mc��EkO��\
�N7b�~3���5FZ�e)�I:u��Sp2'4�
�W�͂Q�B�fFz��7��H+�����¢�����IϪ�M�r"<��r��u�&^<�us9���R���
gƎ���J0��Kǘi��v+�]�.\�orS5�w{!JܹV7ɲF��+��ը̼�?��O�[�Y<R���H(�%jӖVU�/٭Z��K5�"��`��K#�R ��e?>jH �pHj��D`�ܩ�z�Q'�@d��[ذ!´[�zW�2��{�a���y�ב���-����O԰�r�Z�k�\
������y�S�Fo�zz ��i1�G|�;���:���D��+=���Y3���E>�O(,hҐꈼ��^�NרU4�l@��߈��B���5���'H�lZ��P��)ԣ[����_v0�KKV~eI��[Z��\Ǯ���;7��{�0��Q�l�ـ��X�S���쩀�^��ۈ�&I�V�|�X�H/�����4k�����
\"|1{D�F���ƫyr���Q{�������w��#%�}/i�!�{�[��!��D/a��1-���D���5�fa�~A�t�8���u�հ
�8ڱ���^@��ꍠ$�t*f^�38v\A�\�6���T���:��S�YMc��QJ=�.�
	AzYt'��g���dUAh�o	��Y�4:
���@ѻ���8�}�<�eESE�2d|Ѱ�^H��زƱR?�ҎyG��Z���~�Sew �)��|�4c �1l��#�,A���������>+��=���=�]�h�>���a��n@��/�K�Q����#�Y<����`@^��
G1g6�+�����ډ�pe���i����p�W$hn�jM�G7���]���>��2SK��j~��j0>I���,���K�YE�����1RK��<0d֯N�T��5���_ &�jz��.��$t�)����ƴ�e7�y�~ܢ, O��6��=�.��9y�#ē�<�tS�Mз˨>}�