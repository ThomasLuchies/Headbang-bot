��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i8�>Wc�#�?�l��Z�ly��p&zyH?嬏�s��1�ͯ޾�E�6c���"5rR��~Wi����q=n�e7����r�p	��!�S���v�����֣��yATާ��T�Ԑ�s��6O�F���'�+�������o�����x�[��g1�5I�,�R���������M�b��K f%���m|���?+C�_���Ԁ�<6`0(�bU��Gd�$5���P�㔆kI�O�x�� �c���Ҡ��!�v��B��=<�N���X�U�G%h�<����7�ʝ��@�0}��!�v�uHA��^��r���g_:H�'	�z��ò.9��W�@FQ,�04I�o[�@D4�eW,�,B:�]�Ng��A�O�nC���"�^�YK�PM�ǿz-�e�R�_e�O�u�؊l��ꇘ�"�,[�܈B�A,d�v��\ô���-^a�X���Q��d�1mH��-�Oͺ@M�	�Lx>����2�p��
jHT�� �|4���U_2� , ����W<�k2�>1���]��S��`v>��܀�%�D9�Xp��^Z:��bz5�&��V�;�8���(���}$ ' wFl��}Ǘ�qu�C~�x�לX/���9�Bl��(�M��H��<ּ�0&��1��`/�XA��*�
(n�0�(�9N�ѭ�9[�6m=�؍��'�}���zpz|�Sx5�"�e�k�]�)N�$Jpm�����Z�QM�|:�A%�P�%�'���v?�BxG�s_��T�FdA�f4�\;��ЁxoG8	W�`FR��Ԩ�������ӎe׈�f6�9h ���!����W��w�S�ś��I����ag�'sW%��,����9M3}�Ǧ@���NX@ν�J�:�&�[p!��t���א���5_	��,�S7��v�Ļ�Gs��q����O�$
e
��;��&��� ��kܱ��u�����ڜ���q�F�_�ᵺ�#��]������p����Q#k���I,p�D��J,֕I�d ѡ�
G����-�^e�C׹W���
s xظ����tS��]�і�s�w�Z���%$0~ӂ�	�0��s����Mo�Y�(&�D_픐_�v��z��3ɧ�N��㌼�W�k3��J��{v�^:�簑?����[B�e"��6�zm8�>-e�u�dUA�{���-�-���NuU���Q����X�l�ê��ÿ�!�����0�p6Ϩ�,�k�0?�.y1ɔdr8}QTWu���O!�zD�1g�-�-q��3��3�u�%4]�"'�	���O�x���a+vIc@�~�q_4Ui���kc�>��QF�G��Rh��s�#~�����xəxX� �Z�&�9ة���)^�R���N`զ�JN�\�1�E��M��Qc%�]ې�?0ȟ*� ��]�Eޠ����}�9Ae�u�[d��l����oj���?Ci����͓�Yc:{��U����%y�v��~��~lkF*��d��c��V�Ƹ5rc^�W�?Sp�^�7`�Y��ڜtW�My��i�[�=�k(���8���`��"e������܍����0�w�,�q�y�^��W=�D^tb~u���}�jo��������w�s�pi�`�A�o��j>~#ް�E�-u�7wjs�w�a}^����_̫��y|7a߯T�|	ۛk�e܂�4#C��܉�>�Ȑ/��]��<� Ҙ��V ���;4q˔¼{R��]i&�ϢJɄ����i����rX�eR�F��G���?�L�[�Z�N麟�!v��;���h���3H���ؘOU��hJ%5�E����U!�����]��z{P����NgBM���/�t�{�}Xf$�-��>������e�/os�8*p�ޝ�e-��n�p�y��4��N�TQ� ������:WF*@��8���L���MRv~�f�$D�,-�4�p*�S��<���t�|�<��V��,��4��6se��nӤ8{	��R�S`g�+su��%�×T�(#H���v�$?�+=FSpp�	7�ʱ���V���]'$��\7
����g�b"���w������Б��X@� ݸW�/m�r��b��`S��`�:6�.���"�C�b�����mx���["#��,_�)j<�K�*�si������_�=b?q).&��8g<c/�V���؏j����:��f�W�zfA0[+ӛ:���v���
4\�s}�����=�*�]���fUW#�|���v�ƺD�k
5&m���ѐY7A$w� �+2f{����PN��L0�̵c�j󰊈0{G]�кz���)��E�n%J�3�o��[^٘X?���*��j�Z�S��Nn���8`�[Rj�v����$�.��.g4�;�����$�|�r"���� ����b�|]��4�;NP�L��������<���l���3��x��K2dY.ݯ��z\�p/Mw{bt�'٩$<���#���՗+��zț�F%7���3rf���x��?��`p�ר`����!���*����W�%2��.�>�2Մ4xXm��r)I�Uo�cb	j��4�񜦚h}��f9���&F�C��mnjZ�Q�������4�4Hu8K��n��}��|ь�u���q�%�Y�[�U��_�U��:���%�q�`�"�SS�S��|�y��>���˿Q8�K�t��m����~���ϴsxo��.��+/_�o&1�ҘU�|����@��iX�ڂ_p!�.U�ݕ+����%�m�n������<��&���I�ᘌ[f�C���#�,��
�W&+#���cb-���I�����ԳRX~�(�L�b$H͊��Q$Jvz
��o�)�^F$�a+:�jӸ^�7�5�#����<W�w�7�����ӆ?�<=�u��}K����[�,������]hp=oXN�-Xk��u~�?���h'E*��]5����o0�@q�S���a�cC3S�� ��p�	��}{�E��Ԡ�1ln���3�����n��[� �ن)��'%�m���5�j���!�l�E�ո����W��Yp�r}^��f3N���QKP��34w3�����#�i��Li�"�wZ�SYW�z{��5WK�/Mg����{ͳ�KTN?'�CAl;��3^b���i�YB�ȕ:լ�Pu�5q
t��R�ɳO��k4A��?�iS���R�9���zi�4���,_S��t��+��Ζ��3X}z���/���6r�!!���⮞��r��em�ބ	|�\���%N�x���+���=��!z$%(8ڱ���T	��I1,����/<khp]D��������UJC�m��)!��F����bl{B��W�����a^e�B���A��L�L>��|�v>�it�%=�8��^I��u`�vRڣ �<1v�����|.�hO"W]`!}�.�V�p�[���U37��Ό}�P�ꓥ�Mp�k�"]?�b���J�ק2��Փ$��Q+`}Z8�����Rr����1� _SU�cLWG���fn��g��6J�O���U�T8�@�N�r7�D~�r����5>�n1����B����L�֒��ټ{� >&.c��r�y�u�3zg�_:>�}R�F�qst�䏗ǡ����N�g���	o�YN<��~��Ƭ>[�$Y!�z�_t�vE2lJP�����}g�7?�%r�?E}�q0>_E5�o�^	�cT�B�mUL<�dl�����ύ�B#2��M]���/1�l�y�Ƞ��c���Q�@G��t��u��xc��0���p���)��f��t8�C�ɕ�o���0ŁY̒i�V��� �@5Am���;�<��W��7ex1I#�E���,���l0o[[{�.pĝ���.c�JbF� ��[��%�,2Z�>��As�%�3;S�F~1�p�3xTV�bНѴۅ$<i���Ða�(�gM�B�Vk&�r���鄪�:sEfч��s��$�cT߁�'[������b`�ec{���$\W�~YwA�<�S�B�K������H`�ѩO\��E�l ��%G�@.�
s`UrA��~N�o�x���*���2����9Ͽm4�>�ʝ�j
&9�����0�������hx�z��JG%�)HdT�+��� Q���/t?��b1	7��XU��*�fr��hG,G�Z���Z_be��Ϸ���:x�r��꼙��9q�����TUƭE�x��d�G���Ps8��Hs��F�H�`�+BR�5E��>,pl1�xJ�dxD�7�.#������$�XP��h��_���wa��pzK_F�2�x#p%o���Z��q����@�w�$���0�똥kX�uqԢ���%�̤' �o͠��b?�9�,�Q}0&$&������c+�g��K���L��7ՠ�yDRU5<�y]�`͍a�X���J�����gb#r@# �(v�Bm83H~�>�//�	'�x�W��ѫK3j�*B)���|Qf��
[� Pp'����7��u�2�Zc�^�`e]��4L�������=�f޲�p�)$�6l�i��vd�V���H��t���f�\�!��<A���}��S>��X�՟�/�[�O�UvXLv�f��D��*���=� �H��
)�i�8Gy��8T��:�i�k'@��E���z�:�,��<H�
��-qlಔG5j9�Vܿ� 9�$̇�q=B$ho(�41`��F��2;�>�7�j	�(�l�$d� ��]�|t?�k>%��>!߃�A^"Dk��G�K�!�/C�E�z5U��͑j	,Z��&˔��:����ߌ� �{�_���3W]jf��>W]�ӓ�@��g�m����pf׶��V�Rs��P�1�Lpp�� ���!�,���w��q#�5��"�(�}��]G�=
�0H�4��n�LG�w�t?޴�\�|I��.3+l��ك|��s�Vk�%����Zn�S��2ʺPp��g��O��;tO���x��s�z4kX	�������v���ǉ�t�Z�m�%)Ç^��"��_�)G��xGf\��g���ƓPץ�Rij�k�j#gS��,����CiAc����1ά,4a�͓�;$0����]��CV|���y;�z��8�d*���@�N��OT�8��^)�G��A㝌vN�TE�n���P��r��%��HP%u�`J���LP��?�Ң����@K���͹$�f�w�w�n�y�2����P���j�P���!�@��h�&�@�"mP�_URk�H��8d"`�iŋ�N�L�}��+�I��s��'2��%:y~�-QװY��8�;/L���>�B@�w�~)=ɞ(�i�W�!��ܮD�;�V��@g���?����%Bi"ZF+�1,{���Жq��*��x?RO���h9��)�>�������Er�e�ǉ��AH|�r��j��Lc��]�f؉R���.-nO�2�eD���Ì��0���fWޚ,GG���Z��l��{��=U^��>VJ�8SX�qy�Ֆl�&�_�
���Ɍ��2�S��0p��.��l��Z"����Mfq�|�r�Č���4^�h�"�.��o$a'��+ 3&[}��?���e@�z_;��^�C'�-+(�7�4[��kmMd/p�B�F�q�r+F*�4��n���.��L���,��7�����s��z���;��lO�7��Y_�R� ��V�R"8ڙ���>Eq�Ai+�r���C4r���&����:�}x����@E�FJPp��y���{�����v� �c�`@�9 ��>^���F���pE���u�s�Z�o�"�����>+2�?i��6`��S�@�#F��
*E�9�^xp���?j3O��:&�����x�}\�����5�
OE�ޭЏ��Y����� +�޵�C-|K��$f�98\HH��\X=�S9Jm���Ӈ��ݳ�N��4��M�.5��E!)��2"cȔ����yHA��g��ZM�j쭽�W����;���θ��Xs��X�(��A&*�, %R���_π��W���b��O�p���- �9�2d��:�A�^�I��-�A�x�V���D�Q�������'�\��{J�^�\Bpԏ �J�(�Qg��:��Zg���"T�������8"R�$<�Wx��8�t�\ ��#��2tߩ~m�˸�M����0+��@��'f�z$����t�7Ue7��w��XH	�0�kCu3^����O\?�r�f]���:���������,\ԻX�-4�
�O���#�$֡=�J�\%	+Q3��M��g���E[���m���p�Q���G"ʙ �y%�(�X�%�j#&I�{^�)�7�)[.�p3�������t���$L�E\����FcOc�"�K*	�
�{��x?�w���$� D���NкP�P;t!��D58E��iv�W+��l���M�8a�����R,=Ra[/Q��p�HH���^���%U�g([?�\d���e�;$&��D��BCQ�&l�T\��	��)�v�ĜD����\Ctv�k����hOd	R��3����$�LJ���,7ZrT�g��YBK��UO�Q�^�I�ca;�{�q�`S����t>eFI� ���9���2�hM��;ƌ�xϩ$F����`d|���D�n�/�?��Tp��^Q�}U�-��0����fχ�����?�mC͈������2v�M�i�nO}[�50��*P���\1��*\�d�2��g��_"\m�E:��m�֪[ml�����A�.����J��l� �4��~����{�M��9��-	\k���q�i�ԯ)�˅��t�q4 Ì�f��H�6��:�����E��-Y��xKe�@�3�G}p/�Ģ���t���f;�ϩ��(��[>�b����:�)��%j`Ưn��}P����_waLt������I�E8��pv.���Qs`��t
Ak�ĉaR2��`�C�%���V ��4�ħʹpU�JF�;}Ɵ�;��@F����|��
�ya��P�}�h�qdL���`�I��'̀q/X�?�D��J��U�R,=�Ձ�XsU���X�ma0c���e)!S`�Éb��H��87��O��n�	�lp��{��T�����¤N�M���}ٳ6?mk��7AfV6;��|-��c".
��تl�0y_�K��L������!�d~�|�I�gᒩRuD��$Ο��	󽦕�Do��M�TX���3��e�dӖ���쯲������B��O�X�Cg�w�,�,���d��7�F5I���,U�:��VU�B�3F�5"P��d}�\ס��ƭ��K�w���t�����W{Õ�қM&!���b��������c"�������<7O5����vޯs�>?�C:��n���j*�D0�]e >?16g�9J�K��y�I��F��hyB�Y��8gk���*���_*\rz��k��*<H�{�=t��v��_
��A0܎�Y2�"ȍ=��.ue�C&�!U������?d���~�*F���z�׌����C�qf[��I��Zb��&��UG�6�����s[�� ��;���}G�ɰAF�F��9��<?Ѿ��=��� �Q)J�-��]=?y=nrK��~!��?�#WPaz���D�0��^�E>?ʂ4H"D����~-�9�ꔺ6������~D+�@y*�' ���D���;��N����*|.�yʙ3����?��u�lkϓU���9��>G�S��C�V{~�ɬFfBS��ݹ��Y�
�#K�F�ʣl9����J��,��j���Qr�|��p9�}A�#�v�P�1HJ��1��|�T��ՠ|��Nb`�To�K�N����?k�_j�u��2�I���˿m���3��r����-,}�C�aĵ������½�q#d!f`��0S|�=%Hj���O�z�P]q�����ɞb/����߿��MR&���J���@DƔ$Q�"��=׃N
	��j�=n�˂E
���8'T
�2�ʹ���(��tJ��?���=`������P�&c�?�9G����һF�� aU�[n{)?7���䎹��1e�%w�ʸ� Ϝ0;�+�o��[�|в�AwTPu����Z�6��|�^mfi�M9[��u��G�4���d�˛�l��k4z\�ap�E
�km�+�xp��*���lׄQ��GϤ�lX`�����6� C�w��8�J��
�e�sΤQ��0ԿXV� >�O}��q?��".Q���I�3|6��E.̜����)�(#�?�D�ySYY���o"<���3}�!S��W�x*+�S(3M��R$�$�t	D1NZb&-��f �R����D��$Am��dzg�i8��ɪ(�m���q�*��:�u��SӍ��]樥!��	S��F8��b�g=��Ȯ���ɖ��|��I���k�{-u��>ǭ|Z�W��_.�=[ӕ�/�gf1�>�Մ}<|�;��Nmk꣔#�0���_�y�>���;\�� �X^*���9B��  �����l`��'`�\�`���D0�� z���a0ux�p�E�l���*`�z�D�{����l�4溓nA��������S�b�>C�2��ob�(Dr��=�d�cg����x���c���w����UNB����H ��&y���8��e�77_���\rΣ����>V���y��T`��v�@�=�8�k;��I���DߊQ^�L@]�����[�5��?��Q����oZ�.��lˤLI��Vg�(i�w5Vs�00~\�C���(-ǰ#�G��W��B�K	���D x@���'}k���HD�_���,��c�̃j�VY�r��B��C߉����qq!M�3�0Vȏ��%����Ʒg���,өa�JK1��e�-����ld�S��A��\�Ǩa�r����+�\��W�9z�,oM��Nެ�+:<��7��a�$�k|-�%��$K�����b���Ũ���2�(��#��`��z� T��]2!�Qg��ؾ��}󁏡ϫ�[)ȩ{~�w��B�h2��cӿ����.��R�����]��7 �8uȸcV��ia�DjP�3��v�4U5Y��@��-��r�Րy����;C]����\��s�n�  ��s�`�'�<���(+���� ��{���|_�����FO���}�ù���s4A����H8�W=���LO�����	v�)�";��fvm!B<��H0���g���
C�Bo&� ����(���o��t�(U�:�ĳ=Z�\a���6�K[Q�X�b-l:��\)��!yG���'3�<D����@�e�����Փ����������9P��Y�=��1^>����D��v�־����������R_��'��:���7�d߲X�Й������F����� ���ۨ��U�Ȝv�P��b������0}>삨�ź��(Xԙ��B4�������<��%���bn�����qZ�
�-'�F��qצ�-c~U,�(�}V
-��`�>�Ú�jyxGc�����<A�A�h��^�LG�|r����������ȭ6�g��l�&	�-��k�R�v��c�R_ϴ�����O��)3q���`�2(��9����r+B>��d�ƛ�r/;ǡ�A����yd��3�]�ܢ��{�-��\�m-%7���f��#fY�������[/�B����oɏ�
�s	�c� _ҍa����_P. .�Fi�ȆW2½:Ѷ�kLw�¯�x.(�^�"�ʻ\�����D�I󉽴Ѿ�{�E'�hP���1*Y!*�Fh%����e3�϶����]u�M�]-W�	����V� 	�
�b\�Y���Ò���@3�$l
���eW_�OT���e��~DЊ_r�(s�^��R|�hbI�����c�e��E�?�8
�\���:d=M����LE�p�����5���;SJ a?ux�����-�1i�F)�@����s�����׏(b�b��:ED�C���,޻d��B��{��Map�#�"�P����G��� )�W�+�efK�er�9����D�I=��F^ن�v'��{�U��}�uS_5���V���t٨|c|h�t��=ke_xFrFk6͂姇9�u��ƻ���^�$��;���-�韮pz?�"��(�ہ�2sM ��k�A��a�b�.Tc7Q�>f7����SՎ[��  Uv�Z�f�%9J�;�iS�O�)�]^W�;i%	�Kv8R���XeP}���3Ao��z#��T��!;��%n���s�C�����v�Q�t��ú:�$���Y��s�k;����:�a����MCy�
��q��ۚ�RP���{�ۈ�I�y������F��6��Ω#��mE>�q�7p@t�I��M�����Υ��39(r�-��a4�}т���nV���F��"r��]�d�0�j�3�sѨ�\�A}:<���Q>���>�e�Ro���iU�6���z�YxqJwLbH�4 �&fSc(]�?%�%�ߚ/֩?i�y&	-Tܹ��� j8���LTd��)},������#� ;�A<���8?�0��ü�V��_�dW���r9,�����Opa���7�PZ��f��ͩE�_��!�aBnZ��vEҾtQ{Cr��lх�9�o]s�%����)��&Yd/u�$���g͉�k�@X�S��>կ���R�:��;+���m�L���HQ�K0c�W3n��r�zRB����Z�/�R����łia ]�����j�?y|�~��,��Ñ�:ZUt���Eh�W��H�N��*��t�"{X������l͹�P<O�)��*�x?��Ⱦ
���5�w6P��C��,z�F"��y!��iJ�ѐ|��h��׵�s?>�KΚ�#��n�_�u6J��a$4��Ԋ�f�U�[u�:�����?�:Q����i�5���<}ϲ?��{@J܋���N. (���!ņ6�}�|�<������<�\5& �H���1=�&�b��L��I_p���r�J��7�%�֖_���P�5E]���z�-`�H[1bޛ��0'�A��/�ݻqt��c�ħ�K���*Q#�|�I�Ї�	��4n�M��*p�U��~���w9��ꪘ8�M���y�Vp�|皤F��f�{��B4_��-��R%��3�A�ĸ[4��D��a�~<P��FtU8�CK�rg�N�  e��_^�W Z
dK�$js���f�m��q��$���'ː5���{�z����������-�`Y�[M��0Gu	��`�F�`�R�����c�S���x,<?eC�A��|������Rz/ZXz�(수H��`p��G0���4(��H��G7�����UM���1\l�e�a��H�ؿ �]���/�=�4ey��Z=z;@P�Cy�����+1]�g��6p��Ģ�v�g��t�Nj���ת�ެ2�I����<CvT1�mV<�-�}��@%�Ng�"'�<���[�˪s9K��34h8�$˻�l�Zf�h=!��mBHG}��;�9#�>0����;�|��5�����:QeB�h+B���L�7zE���"/�}y�|������))�Y��<�o�Y(3����o�c�ܓ$G��R��4��o�WZ�#���1�2,���߷�]��^f/���	25�Уq���-aF�`"&�}��gu:�����9�|P��ƵB2���� �}�*�p�c�o����6v�O\�`��/����r�
σY�Xq��Sc�O<�7w��������|�|�s�P�EN�
�s��@�e
$���X}�V�g]��+�c����������F<]�C �cE'�g�-lk�Ek�1ܥ,�CX[�!A�φ	K���q��8��o��=�:x�������Xl�b8�p<{��8'yuw>N�sPfm�ʕ����_��$��'�!�q,r�F���& �:��k:uʯőz��K:������I�$m�����uGP�|�a�ns�u'+T��Ds�a��G�:����-3O���� y�pٴ&z��J_�2���~pv�4�[p�ʽ������.՜���VW�5���]
�/��#p<�6�<#�,��f��P�LG�1b���V��*ʎ�˜�3����F��=�\�6申q���Q��1p!�E��x����(۸ns�~���&7}>C�Id�}�I!�ٖ�KJ̪���{��A�a��z㱫���$��D._w����,�9�u���#�E�>��qd'���7��3V�4�h�[���doU�ږ�`�J��}\fۇ�Rv���P�U%��D�Cwy2�3��+��`��1�q���������j��>�=�j+����
��4|����� 73�4
����$�,�Ryja`c��t�Kُ����1Y�?�'��w��m�c�'�~@��q�$2�r�|n;�`@w���(A8z4M. �A^�wT�a�_�Q4�½���w�ڎf��X=^��32��a��ǧ��{�N�B�GILd��ځ�9���F�-�����N`6��n��>6)�),�=԰*�u�KNBC<^<�1m ��jE~�������Z�N�F<n)�PW�ղ�u�,����̼�?�v_���#�(�=4.�:k;fXs��:1�Fy��h��S��|�n�N�,l�Ż�}���wA��v����3�|�������@48�������S)�������fl�"KԲ�˷ob7�s.�c��Z97ts�3ۢh�ȁ�7��7�����=���+�%E:3�����A�iG�A^2aQwu��'�xX�\����SB&�HNy`x^���何��y;v�\�y��7-���E�U�I!�"���6������
d�&>�n	DswgJb��:���tg�����[��D�=��-S��P@ ��)�2&\��<�1�=��W�>�v��)7\2re9ͣ%�#Q{a-�m?��B��8D`$�M����5��fDA�Z�nX�)U"wHе�-���ػ �!SlLN����
���nK]��I��P������C&p�C��e�����W![)�
o�P�aTb��Xu+ن�"�W���LAm(Dm�����JS#A�@�#�!�ו,f?��� &)_�j	�P��!+�Ъ�����A��Q�`Ⱥf�l40�=�'"���`Tz��F��$��[�;Y��a �_Z�X�>�0�9oS����ה�W�f�d�?������1Y��{��q� �v���{Z��[@7�&s�U� �N�f#LS
Y[�?�ēѩ��{<���f�;8��3���eG�e�(eH�i�L����(
9C�\|L�q�kw�o�	��f@�Wg_v��N�(�%ŅN�Zع��9�^*�B��r���4�U{վ*x����(��
t��B�C�S6F�ͪm�X�*�3��Ǜ�UOy~"\[ࠥ/�u���s��)(K��g%Ǜ�m��ۿ_?~)g/�{�Lc����#�*�ڇ!YccЋ5�x	_�{��r/6(_b��Ҡ���ܰ�%%@w�.�wA>gADK�ÝV�vG�����\x`h��nv���&vRi�{�MxUZ�˘k"`pzn����n�階P��hհ��r�`59���7b�]�?0ND��1��`���l��ϑG�3)<���҇ 9u�a�]�M�e~�Etl��rj� s]��g���4jJPQU��_������Jk�9.���Ԓ�ǧ�T�^S���[�O�,�u-�s2�\{O�/��`�q
��KAc���NyIm8������k���fu��}�bQ��ʢ߂ˮ�RSѕ�c��б��i�5�k?Gӆ� �9w8��/N�T��(��V=,�����]��˲BhJ�R������# I��0�0��h�B��]�#�'\a,Sl�"��n6�N�Y�����W?{���N��XJtR�� �CZV�x�_��Z�����+�I�:X�yrPX3�8�,:�����%�7�M�Y��cZC������ �y�_(��~��Q�7�1T3L��轍Ɏ����qEw�
���c(I u����d`�È;3�'�9��㐍h�s��)2��[�W�vc|����rQHr���-@�L���X={�k�cx�8FA컬y������|,��J�G��@	�l����	Ave y��9(r��/5�|.Ә����7��i8��|`���#f���2C�Z��,���М�w)�ΑF�,3�h��!z��U��q�Y_�w���t&��LÇ�� �I�0�x�J�{:���L��g����}�_g7t����&2�
Lm/�ｕ�Y����{�#��ők�؊9:t�����giM�oQL]W�y���M][ц�ɟ�$�S��Vƚa���E8��"缟�7��ٶ)�S��I�@�������:�X�0���!782UY�~޹Fn7�z�3��HJn/�';��Z����f�ff�z	�p:D�z�{eǾc]Ƕ�RL`�~r�C��Z��yz���=N��V塞�\&t���u@�' �����t���
���	/�(�U)��o��HbGp8:����Ny��L]���W$�h�����Xqk���*ӿ�-�O����Tldn���6<��U>^�N\�I����6W�L�kmV�D���r���W�eʎ��b�Pz�<CGs�􌢂r_l�|š�0N,~e��dZ��N�b5���{H���g��&�ֹ}f�y	��/�2�Ӡ�W%m�������s��L��*9u��ӭ�S���)����-a�!�'�f�+ywg_i�@5�B��2�ʷ�;C�9Q��ȏ~�?˨�� W��+�9�_l�M�����y~�������܏ �x+�Щ�P���3��״ص��$r4�X�� zLB���͡�\쟫�	�����LkY���8��0��?I��&L\�ɰ����sГbJ���f[(�BC��*�]F��CK�I�?���^5
�rui�_��fgeMl	|@t��_����������K�U����A�'c���-���R��O\�Y�w�R��f�G�AqM�$^J�U(q��4���.�+-��y �U��$��L�G�F7�/�ۮb�[�$��Oх��a�iW��R` ���9i�.�,j8���J�fW
RS�ה*��.���Et"�X������6��D-7M�/"�<K�/>�O��e�}бl�|WOT�h���?����Y�p�E��\���&�!����|��v�.T�f���ɼ3��[�~2��2mG��n�r`I��,�%T���?1�E�~�(wʕ;�����хo��P�í�"$�{8�c�a�6���V"M&�0i����v���[�p1D����ԿގiI�o�b�}<eߩs;e��(�'�X�e�e��eOLH&�]Za�,
 і���#P�97�=��#!�Ԣ	F�f~�f٩&�����0 �H��H"�