��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k����W�z�N��VXi^�p���d������֡u�Y�"�׉�.:���O��2K���r{Lٝ���1f���^P2�8��ۅo
�W4��6 >�'���ufR N_-�f���w�B�t�"ʪ]��p����@0��%�\�$BP)�3�H�ۉ�R�y&�w	ʿs��� 	�Cb�{�_��k�֦��䜯B�[����`g�����޹�v�h�[���{HwZȔ�X�JU��h,�+�Eۋ9�5~<)6�[���,��;�2��`4����Ksp!HUN�7j(� $�4��R�鬤��Noe��.5��zN�_z�(�i�X�MQ��'4F/�U�g�F_��:`Oח���PwS�����	PQ�#p�������O�M3/G��j���^���7[�cR$^����أ�N۹��K���u��Ud÷~/���-`���h�xŰ�Q,Ќ���/�0��]�����xW}p��D��O�T.�)E@`2�V��O����f�QlfB������)�(l%z>���.yR��tD{����~�c���=���+m|D�^N'8\�'�=r�%����;�Z���vya��v���f�i9[ձ7�^`]���L��y9���������<��H2�G�w=f����V5��~b�W
$����EXs���ۂZM�8)�7qR�;B�0���
]IN��}�!C:F��J� d�y�j��i��� *0*'�HM!�<�t��:T�!ǥ?�7���K�\H��[�i��BR�O�V�A炸�U���ex��籟=�t�J�� �w�<5����(��v�}��i-%@ޣk1���"5�R�=(�]��s����)�k���2�f�7b�W�t@y�{�"`}?���֋?�j{���f5�W��d��8?��m�LO��G�h~�(cٙe�� �^���}焳�����,��8�)�a2��/Ֆ@#X��=�lnf���z8�E�V�]<
��������UH���MH�^�y��B��p�q I��i��h��薑˜��5I�u���LÂI�w�@1�׋E�uptb���W���m�՝��D�/+ �Χ|�Na:�*s�[���b���ɛU�?=��oF�Ɇ%�j;a��O�u�������:�1�y��`��v�|Ē�=�_�&J�����������^[���Wg���_�l�����3� �K�<���),h�~%Gˮ1��x���?��� !� �/����s�pGa.g��e���H����-MA�0^[���.����զ3�g����~�˅��+�M����_ӿ���V��+�v�K���>'`��ʗ�v�
����OJ�(��K\�ꒉ])ۚ��4R/yD%����Ѹ�a�| P��� �C4Qifds�껸��`5N�@�)�"���":�/i��`ۀ_�?�U�3G�����_�~�s�ת���Y�����y3�w"�'A��N�f�/KIx|�Um~��
��TU��Y�	`�߲���V�kZD���q���ǂ�qp2�XB��@��R�El���i�4%ӆb����,U($F0��Bh�\{C(�Sœ�j�B�<d�����c��%U����)��-Q�Vҕ�N���kE?����$5o�Q�|�����7�pEsK����?�����S3���±��j�צ�WKq�����[�h���|��#^��19���)-�u'̈�7�,KD]
���4}��	�SKM�iݜ%�f�SXX,�DlV�9>G���s��RS�����O:6*��"����uX��0`辎�����&���FS���e�=�ް�%R�no,ݠ*�0$$`�N���;�'��\Mߺ��/ ו�U��|!V�2�H��������'� ��F�|�'���&x�wZ�"�_�2`,|-1K
����%�݊L��M��4d�[�Fx)�[�0#�tr��A��z�\�]f�Lϊ4��Mm��I+l���l�yI�*,�D�x 3vި����E���3gM��a�,F	��F䱢��A����P۵�n(�4� ��l�w��>k�.���+y\@���㎇�'κ5��H��Ǐ����%���Q��%q���O,#*���|*J��w��(ߓ��P�'�,�"�~s��i�vS�Xo ��8�NT��o�"�*�.I��Df@�D�����B�;+`���\�ľ�1W�!��΅^���oO�E ��\���g�_G!�/u�'�i�>|!�Nm�b##�>�ct[�vw`���v]��k=($-�����aJ*��Tt��1�kV�S��i*�w ���]�]�
���~�qkS�3I�% �{��J�Ӎ��+�w6�N�b+)��V��
f�\��3�|u�X�dJ�qN)�V�=�'��x�s�y���u?��*�ĂC�����ŰHB�Ê>EP�đZ�P����%�"�ƝF�It���M�(�>���ҊR ��fl����ő�|�B.��#]�f:&8��;p�
th$�x�EL��>����PJc��R!�K' �k�]�������� ������w�O��/ӱ|h�
p�������F�l5AÇe��T.���Y�yj��<�����eI�
�g�g�ܸ��)�-J���]�sW�o,�K#ߕ�g�����IF��В�P$qq��'f�K��jF�N,I�]�nFb�j0h�;���_.T��-���C�6/�3�P��/���Y�jǫ��D���I�gVɂx
fy>:O�j.�_"�#�c�x����K>�J?e����g��#���L��3�HJ#�&�\�je��������Uh��]��/��ӫ.�K�]m�:E^`�+��������B-4���~w�3.j����Ծ�����H�i}�-�z�'d�8�~3���;%+��6~o�^�PPS�fS���I�!���Ъ{G��G��]tV��}1/��{���|��0bNl�uD.�J����Q��Aq����l��T�R�'��B���;`�P<rs�Ӓ%L�����%���߲�7ޜ`�@���;���k�g�x|���'������}� �W���hÞ� �@W���(j9Y��!�~ik����X㖠XK���.wY�4��h[���3�6��3O!���^�����R��3�H@�='Z�dߨ��T�۞�3����p���AG[��nE�V	"[d��H�0!`�6 �K.f���4]8�W�ؔ��H�=���!�^���{�pӺhȃ5!�s��](�(.�ힿ�@*���pb?�Z�E8�����|�!�ͬ�L��7]�` /�
Y��
��p�9�9׎l�(��k&��6��[o�S�5CE[U{u���h때{�y�Ki,���X&*��_��B�T`*#Af��=�ǨH;��7)�[�c���� 4�j��ӛ��	nqhK�+��;1_2F
10����֓u�c�MHBo�쿝�Z�u���\�laUծ*�6�����u�!�����Z�uJ�{�Ao�!q�Q��Gd��� GUq㓍^�YD�I���Z8�Kx ���˥J<��J���"� ,Ԁ"9gv���G�E�j��;�f�@10�YM�א��j�`��T��ӕ@t�&�� <j �YMX��M4��{	� �-�8�Abs�>� �h����:�t����G��:�^���>����)Շ�E�J�C�Z�Kli�vXtC~	�ɖ+�9�v>d��.G�OiՄ���L �%T؛'�[��I�.�����2"^X?��_y�:�E��p�r]�P��Y;�.���V=�!`��P��D�xR�i��L��m)+����RBYCDt���ZP��<�f��ۨI
��b��)1n{}&!��/�-��E1$OO�y+��wn.�>2�6 sR�;�&�k%A:r0�MLԅ�{%N[k#j
S: �1/��L�C�aOǦ;uG���XE�����C��G��%J�U�R�|�@4J�H�i��*q�Y�;�i?Ơ�J#Zs�e^��d��,8��ONϭ���ݳ��c����U��A���ֱ�o���&HxYl�ݬ��J�-�5�B�b�`A���5.���	�
�޾x޼$���s��eI��~@!��a��s��ʰ�x"m�Y��a�H���ѿ��}'-���v�U�	c[��2tI��L�����l1����/b�bx���5V(fq��+���g�RR/��_bQ�c^��9-@�S���qV��6M�5�-���	�z�p_�$#�&4O��rT犿-N[��Mkw�"�4���B�����ǍIγ���<'n[�t�tAg����J5�X����1^���k4��&g]��.���$5�I�^(!'�3�"�ԑsއ[%nbI9R���]#����]�*,t�1�<�/��M�|9�o�t��n�6�s�9�C�������`6p7b���Ts/L-&��Y�Z�� '|Uz�ɞ�s+��hD�v�Nr�?�p�C(���Zy��6��5�)fwlp��:ܭi�t��A��TIU�Q�tQ����D*�p�Z��r�d�KG{�IEq�� ����/�]~4�4L��"X�xe@���W:�� �e`_��T��q�b����$�Q�:�bn	T�nO��ӜW
����n����W���MWx�p�7;��_g2��N��%�[?��w��(J�&Wb��z����;B�w�h�D�d(�?A���t1L�פ�9�m"6��x�]C�����^�G?�1[m�v�9FD�=7�P�:�?��� 2�[��wޚ�/%��)�ӷ�w��N�o���Ar�ܳK)4VQ���M�?����F�b���(�D&�t�#���H�C��6�!L"��XB�wȯR/��9�q�5E���{0�h%kkh�S����6j���hiU:]���u�X�8m2�>�aW�qA?`��oG3ʡ��[iU㤿n���yϻO���@�$<ч˻ V2�����,$=`�~a�S��򿴙����tl�C�ju�g9�%
)\��?�ށʫ%���|c���L��D��16G8�zN���-�r�&2;��	E�/���.b�����t0$��Pǜ����+W^�ԿB�vbC�ڨH7�*0�ǳ�}j���|����P�"��	���ɻ�~����5�*7n�>��ݻ��C�@Ƭ'�ԅ�ԗ5��3��G�N��������Y{sIQ5��N�ِ���Jyj�h-@|v��ޭ�U�뛝m�so5v�:�h�(N�ː�s� �'7�Qxϧ�5D.�|Rn�Rl1F�-�tA���K�u�$*�:֟��Sܺ����ۛ�i�qI� mY�b���-��X��"���������Þr��k&w�����1_g+Ly����k2�3��
��[ ��	����1ǣ�%&m�VаGh��zt���V��#f�Ʋ�R�.Z�����s�Wih|<��a��� 0��I+�Y�l�m�Oj]��J��"ȁ9�NZ��(([�e����M�oC��(E6O7�T�]��qK�3J��305S�H�7�6��ۍ�eb"o6]1�B>s�Ҥ�&���=��cHi�� *b�OAN�e�ۨ/���YS�8�-��g��0Mk������A��iү4��rb�N�v<^|6�|Vf	�˖P��b�bq�����ڹ���͋�E�:N�\��UU�;,q�f*��4K�t�����k�>a#�"6j$�J��������RN��v����r�MA�߸!��h��1��nr�
Ht��{U��b���%*ļ���n���x�Ļ��L�)i�32���.Nv��S�Z J��_.����T!�"ry�}W%��-� ar���Z���aR(��$\��6�\��&l�G1�V���%����W���곜5i���E��H����j��;~�3���W}+�]��^����������u��M�:�,���Iz����|�
M�N��Qb;�c`��`�G�o���e+�P`���S<�������[e]i6�J��l�{���P������A��-͓�VB�+���Z_���������	�]d[��Wo���)|�S��x��(8JY[�I��Q���7|�_n�ĩ!�6�ˬWCՏ�GZ9��Y$-H���U����/qqD�32���5��
I ���|��g��0]�!o=EK�o������*�P`��:�����<3mU|s�S��:"=3J�X��^�OkÈA)���+���L�q&�{��=&��Ca,al���`L0��v����p27�����b�0�F!�TT���6;z($�8��Ӝ�#Ϭ R{GL���|�d`c�`'�|�l��;W�Cn/�L��A*?N����w��4��U:��h �l/	A�0/��ؿS@�s�V5+t%��O�F"y�<�9|צ�Z����
�\&+u�!�DE:?��}9*��0�$�r���y��w�쥀��z��Eu����H��X0PB(�f�Δ�6��3���^���iڿJ�5|����CjNx����g��hR�a�[ � @���#{ ��(Rڿ�6s�N�Ww��bc��eS%�&��]������s*~z:���C�Dُ�=�� '����,tޢa^s�9c��U�v3�&�h�V"�H��)��H1//��I�Y3V�'l�G����a�i:��4�M����Jϳ�����'��9��\���1�"�C�ʣJSlmGg#��><k���p������2@��K����8.��ȃ�)���A/�'�M�݅��Ka�U-�\Tɼ~T�Y�*v�C�a�7���#���qj����B@�L�b�^T�uH�1%�~g��	�G��d44��r/�찖��t�{�������я�u,�@���5Cnx�ێ�����{��<��m�W(I��+���i"U�8m8к���Jot�΋���.�L��g�pT�5C_�+�wL��l�a|��`u���}�ny9�X��Ӻ�:S2����;H�󖠦&Ϸ��xBp� u�ۻ���ͣ��-mzS�0��$�އ�dcO��vq�jV�
��@rfz�j��C���uC�G隕`�[���ۑH�2&#{V�-�܉�]��WS-���J�m��=Ɯ#�Hd��.�#����w��\A|,�{��@ |��gdr���H��
i9�}3htJFp%7��,N�_���4{�B��R�S]>\�BxZ̡����q�y�ӝ�B�W��Tq2ת0@5�ӝ;%m!ʃ�]�F5q�t+ȡ���|�rmLV/�ϝ�x��B��X�w�x�J�EevRpbD�D5y�WG`d�L��|k�;JǲNQ����q0W��w���Zǀ�ɷ��{v�3�����G���7�o; @6�)= ���Z�c:��M�D�� F�u0��s�#���2r�̺�7����hB�d�6�~(%`^1�9�����o�jD�A�4���z��hԆg~m��~��V^o�?��5��Ԇ���V��Z���S1�ǳ���a��4�א� T�"�(��)~��5�
��T�2�R��N�J�+&�D�Q75Y3�s�e	)4��!�|Ζ���T�Z�F� ���d���F;Kos�T��c?$:'��ۦ�Y$
�a�="e��5kVU��9�P@k�9���O��%q�|���SV]�}ѩ�M0��M%xW^$B�J��V��F/�Y��&������%�����)A!�ũD�;�/\&��Uב��~{�y�e�B��(�jC?#��>.��I���_3��/1
fy��R5_G��9/H
5��0|� �Y���%�U������BE*>-�[�]$r�,�Қ�;��E�5���A\,N��|��s��a ��o;��ϩHJ����*@=5��7O3�PJ֠�ؙU���|r��7�Bu�r?�X������q�a O3���n5��W�������T����:>|��ᅳ(�t�8��&߬<0P˶ �A����X@�Y��Y�4��᡿�V���n���װ����N�O�Tʔ��U�̞b���a����7Uz\#ªOW��3�e?�E��Bj	��=4TRB�}���^^J���-գ�,S�t)��0�P���������U#�i���q�X��AfYX��G��o�WX���o5���f���W�$+ٷ�*�?�y����Y@�����Z��U�םlm����~����^zI��*��!�j5��&���,u��ٲ����:,��t6��O�\�4����|���Cv�/��/��&�l	g]�G"����o�*%�l������(��_�Sk�#.pl,s����)d��'�`uS��?�z���o$�DI�g���{�B��R��v�-wm��t��'m�֫�WH���b�����C��>_���s{v�S�c��E=���1���d65�NI�^� Z���L��0������!3*��YG[oO�����uP��#3�5����X�<���?]�0�_(��N"j��2�8&�����"1�_o�tq�=�K{]�]�zX�����vH����G9�fZ]��w,��鋎�=��l�듖�It51��n�DD*#~�ʑ�Ȱ޾k���o�B-���t�zAH����"ߪ
q����]�H�k��y�Jf%Y���7�f�S/z�/$�r�����:����g�o����{�嚬W�U�it���~ZAT<�g؝W�煟F$
�F������D���Y�BO�+N-ǜ���)�3wM��o��|4�]r,��3�U<��2�u���
~��1�1�
1��|Q�1���	���;��$�3e�U�*Fˍ�AKU&y��;i�6�uL&�kf�(��)}eA�L�Y��piM5��5��A?b����3�@X�JI����L�1�`o��� ����}�1^�H��WQx9}m
���&Skʢ��d4mܥ#���@ike�V�Z��P��`�Ls�ԇ(� �?n�n�˿t���7	�z�aXK=�X
&
�\u+�x�zk1��p0T^ �ol5eml;��*P�z�ؗ�|�1�fҧL���\?�6uґ/��·��ReκG��	�#�1�C�sV?��,WO��;CxF�e7�馃����'��ۧes��zw&ϫ����KKο����y5)��������#����h?S��0�:�׃��r]���A��7�{�����
��Q�gM��2Е�bϳ�.?�^�h��Y���Q	� rS�	�%��Eޫ<�M&�;�8d�ɮ��a�ٿ0`�u~!��Y�ZU���w��kʇ�	� �9��o��J~�)v��C�� �3K}ؘ	mg��7P��3��R��R,0&a���
w7JcD����i�H��1��e|��V����v՗��E,i粃���$������Uy�-ƾ��zk%JR��(�6��@D�b��x�0� 5�t���ʛ�߱�����.|�z.ᡏa]���8�g)��긣{����7��$�U+��s~k'v�j�⋍�F+������Kd��^�L8�s�Z�3)�kL��E�!��k���7�%%a�CI\wF�m�!fB��2��MxMO�|����59�:s��l	�e>A���`�d,�8n�2�G�Jvt��g����/����`��v���������ߟrWķ�f}����)�1�&�~Y�Z^i�_T���R1�y�(t�xiy�wQ�Q��L����x#�l?�2��%�^C��P[	c�O��8���m��Ц�Σ�-������ה/�뺍v����g���ۨ�_�P�����*(��HPo�����T�q�,�)j��Vl��(�w�3,��FF�����v�ڔ$�eT���E扳�#��J02%����oA�+��#s�{*sa>rAV���5/1����k�R�^Rp�Ϟ�pZ�8_1�}�b��p)8}!����ùX��\,���Ȉ���pIe �X6���*�珹.J��l�v9�� ���R�{h����I�@�/�ӏ[w���	�r�Έ+,�Hj�YgH  �t�^T�q��uKx�N���-�ޥ��	Xp�DB#GÆ�l�^���\T����I�bۍ)ۼܽ�<m�Xz�>�O�o�J���?�*�	gr:���>qC��
��2CH{�IH��9��ji�N_��]ԙۡ�<A���<,�& D`A�El��ԣ�lq���E��ߝ��e7C��>ʤrׁ�6�7B�->��� �ޜ�?�8ߔ�`���o�V���;X�F�3tì^���3O[���'��gõ�S���E�We�L�����ؿ��[�4� H��2qsa�K)D�U�잞�c���_��V���M'��Ծ\+?��(�b���°;/�&��0~��3#��y0��-z��@�i[�hr�V������C�����5z`e�i�T��ۖГͰ�r���E�	�����/"���ѓ^j�aC�Tk �K�N#@a�"�P�