��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k����W�z�N��VXi^�p���d���"�f�F�7t.�!�-�p����F7kv����A����r|or�b��@9I�_|'��B�΁��JHZ��(Z��Q�4�3�}czE2'�����e[��$��6��u�i�BKx@.t7"��2��q`��i� ��x�P��D����g泫�b�UVEo���S� �K����ǤX)�w�ԙ�����x���(qx  �O;X��O��&Y78{X1�K�4��]dc����+m+�$��d�$�AH����`LACQ���r��߆7���[x����T��3�L�븮�X���o�7��Wr#�Rט��8����O���=�������x��7�*/���wc�չ=��i�V�V(�~�#n8�눠��n��5��}Z�jY�2~䛷XO�x\�->N���ј]dT���e5R^��=�F+#G
,s�;�ݣE�gzC��M�4����2�v��]B?,�$��%�o
�1nU�Buc�|	a�Jƌߡ�Id�4xM�����ט���K�7f�ε�ԍ�����k%#�o�o�f%U�	Atg��ֱ���<[�����aY���:i�&��i�G2PV��n�[Z���U��|�>:>��S�3ߣ]��V���EN���&_��Z�	6ƞ�j.:hY��`�e
�Y��R�� }q%7:q)��u���L��� �Wd�\Q�@AL����;8�nV���3��2D2z �sT/�K�'xzz�-���)��� �ˏ*C��P�a���~��8�]��qb�h�&�j4G𩽲Y��>6P�\��j�>����=TI���^ݳB���ÇfG_���^�J6���g�j+��� �m��pʙ*��[���^��D�i+\���2��~��mrT���/����G��H(���*�Q�}F��k ��7��{D[�OO�����=�z��<' V����9B׭`���Y�����(���~�] ĳ�3�n��)RN�aR��(�[0H��j&w>�����?�3�G>��വ?-�uJ y�.������./ Us��]_��Ҡ��xqy;[)yHxj2����\׌���U3�:���Ji��]� �rG���z�eQ��m�� �ˬش����%�K�哴g�L�ݜ.e�v��y��]�\�_���逺����X�����D�w.�س��Mr���,�7�̽��lߜY���L�^����1���2����a�P0��߄ĺ�.��
� �u���r$���#{�cG"ꆤ���zSy�}D����>���}+ni[���!����P4d]A�!�As��y$��N���jL3�x7?�}cot��fxc�]�<'@O�X�!⁀X!F�F>M�2ܾ2=b*9s~a/kT�Ѵt�&g�N[]C� Â��]K�{P�r�e��^zQ�0\�����ɢ5��)�r�Ө�D��F��x%+1�KA�[��|��]@���sU�n�M_��N(r\��+1���>_$!�f1��S�~#��]����#J5F�4h�Ch�e��Q��Vm�?9В���-v7(���9;�G����^~�8�̚F���s�M�B��䤎�os?iy�-X��HhP�-1��z�n��ԟ}�1�t��ͭj�wn�e���6���jz%.R����5�?S���;,y��%��}��5<�����!����E��5	��q�e\>R��F�����v(�*�d��Ϻҟ��GH�ᒣ��$���J��h.�j(�,����ó#���RAR�FK�W����v�og�y�A�ِ��	����G��:b$,��;�*N�*-���Ү�y�&��b�`m�7
��p%*+��D*�n�![��MM���&Evp�'{F��W��^T�_�f��/�P���"��DP�7��je
�}7Y�ot����m ��$�,r��F�ȉ��5��+�ƁS}�z�#����MR�0I�s�q.tte{=����T!�zj�n����I��bC�,r��o��e|���ft�V.VFk=YS�k\�aM�0vO�3;�r2�n��c(s����qA��R��?G��IA�m��l!3�n�+"t�*�oN��Ҿ�����+Ωx�Aջ��ϸZ�U��\H�=u4��PTﶁ)��C����%/3_#�{3.��p��m���_м�i�թRO0�8��#�0�`��� ]��Q�����u����U�B˕�/z�W/X�.m���F�ZW�{��1�S1\* ��mA:4\T?��p����5�g>���U���=I�ٕhJܰK��wK���U2 e�Ճ� ��4�%�Dk�L3ъ��ɒ'�ʘ���.n��T|E�6n�k-W�T�Z?/FEc��p��`"vؿ�P]��8��L2�K���?�aGQ���E����^���� ���NQ��,=�3�/x��j���04��9�d*K%��AkX_<��e���~-��w\���Hi5c���2d�]es�q�\���{������v�ct��hd��a)��^��d������.?�vִEC�h~���}��%j�pi�L��ԝ��:�"%'M��dY�J6�ɜӦ�������1D��G�4��*��@��5���WR�Hā���L��t��u��M2 �P��F[�HA<*,��4sz%l�����h@����i4Z3�1-,d��Ԍ�#����񹲚\m�+�����AٽR��DhߎM��N�1�H��]����w���*����= Jp��=�xH�L���^T�m�lH�WKI������ǲ�}��Œ�M��= �����}	�yʂx6��슟�gN��6�P� 2�7=�����փ��3�9M�v���'M4�����=r�0�K��e�F���y�Q�{t'{���am�邁�)��3"U�0�ʄ@I���@�r�X�={�8�stdE�ҭz�#?�ڄ��Q$fe�xYtG��R�L��)�m����C��`�d�E"�1;�c�O�[E4�r�D��A	���U�#�E�=h�a�>O����]�Ɣ�Q(HqW�&��D��ʎj�}�y��0k��ǌ�x}źd/pr"�s�m�����ۨټ!*�c���l���,mzNM���%D��6%����%�F��m��,�CM���??�I��r�r��\gs�������WPbĢ5z�[��.x�V�	q�1�1�C�R�-���OwbZ��j3p�LT�A=F� ��k���
��Y���J0*�ҏ��M6"���,l���|�+r�XY�,P^fF��H�Ԓ�J�dBf܆���A+��ἪK��S~�$x>�Q�l-a��x�H=�����^*�p�N���3�����T��:,�$1g�z�s�}�o�qjk����xLr��j�A�kVj���9"��U��舦z2�����hR/ekO���b�`}SưߦT�iL!45��W�j�0Y�n5���8�zUN��	��p��h�SH���4ȸ��}�W��!er���j��c	��dY,͆�+�ՓG���i�o(�:�;;��,������=���C�^���(�U_�/��Oy/2��*q��hJݶ}�vB)��%�g��4.HJe�d�jyE�
yH%G]7ҩIR�A�PL=-�&ز����{��j�Ǥ7ful�YzR�v��U4��;����	H�D1L�]�9�,s)�p�]B�wѼc	��������$�>�1I���5�;�¨���O�O����T"�_��B��$bBޖ�x��e��(��u�1HP�{��s��؀о�s�"��t|��NY�`�P������xP�c�U^*4�t��g���mQD��6J���k���(��)����9)0�>�> �Zu�[���ٝ���(�2��6�o���zD��n�F���mD���xlZ}iU�B��!E����Ĳ\��6%@B��)J��p���������o�9ˆ�����d{I�,t��&:��,�z �$6�!	�KC+�� �A��=�D�O��:!��S8;Esʧ0����	���hs��ÿ��
�t<p㻼(���H�}LJq${��s�#�f��\T�ʉ�ޑO��w0��a��/ 5�1�}�So���j�1�꿃�a�H���Da���	� kGɱ��;�a����[��!�����X����Fׯ��N��Z1m�HX|��S:�]����3�gB�n����EQ�F���%
V��ϼ܇�`�2�)�W'5i�V�N�M{�vx�c~D#���	�+:F'�Ps�"@ަ�L�W�l�-j����
��M��K�w�;x�rȠ,�v�0�n�yl˜讬z)��k���!I(���+l�"gH�R�=zĦO'�*������-}�݄d'`K��H �%��^n�V��m*� �\-�\�s-\��-*}�����&�������'���E�B7����飷�X-�&a"G���a�&ޮ�	{/!uWJ}���{�s������"��Pmr�b|~�V�8�n��	��s���sóǾ�e�Q�ۆ���GS+4��Ys�^B�&^v��{xuz�7)��y%*;�t��5�a1���('L��`~~�
`V�o��J�y��u[�c�
悠��V��p;s%Lڨh��o�h,�Ɖ��<l���CYx�h�����%<��ht�p*�_�u��n^��o����tr�͝�լ�K|�(>)3$�A:G�/XS�ßn�ҷ�l��Y�=�TxT���ba�f��'���J�|u������p��2��F�V�2�3T�v̪H.����V��O1h�>(�"KE��ws���S���Yk�ۍ1qQs_d�6��,�/T�^��������K�{t����-�d���i��$K�˴�Rx%�:�P�<�e,O�#�k0�dN����g�^ل�����h6p�3�o~ӳ�u=�ۤ ǌM��������I]v\���74�7%ysc�&�Z+Ck
MW)��W�m�)�]�?p<��w�V�})J���z���@�MGC&������z����ѮJr`z�%�G��~�?ebL�)F#݋N1В�H�F35aೆ�k���p�27�sa;���b�:"���rB%���3���Ii�Nt6֪�A��k���s�'�v���(h�2!�K��<Q A�㌟ʻY����5V��H�K �HA�@�f
��[%��=d��Ar�0��&�.M�,��,n�f	ۇ��i��-k��x��`h�χ�G\�Y��!�<� k�͂x�����F��,`��N��E�Ok"��ÒD��8@�P#M";�7P���3І1]��6,��c�$��d��l�;D�b���_t�x������������]3�ќ�G�����+��;@�Hz{ ��5��]XO^�F��8emh.2���|0�i�KL�
��ߴ[i�JV��T,?yoiv%�cC�:�M��1NW\���zƧ �mj+|��]Tp
;a�~��tKڝ &zHūI$�1����M�ai) j��]�`޿*�/Ѻt=o�8��GY&B�VT��G�}���v��E�߉�?iA96f��A��>[�}?b�Lu�C�	;9�m2��=�x��h`w�|@�֌��jߥy1�pZBA$]�_�m��_R ߛq��������#Nku
�Hk{��d�l�w+
f|W?z?q$�aOK��̍^+ٟq �Ei2u��M���I�|s�9I��� ?E�g�0�����׫v��5S��5ɋ��^���L]���q���sV�Z��'�K�1),�g4\"n�'�p�x��xЮ���.����Ä�A���jT����6:�6w+�fD"t#3���"6'��)�η��f�E����h��'�����ކ�@|�ϵd��#XDf��t��ޑh�G%V3�n ��ʝ-���Lj�az<^�hU?�a\�(ގRV����m	��d�ݠjx��U�\�?��%��Z�`եd���78;���j���B�N�Z���W㬢J�[2�B������Aˬ�U�x�ByA���tUbG�Zdm�Z0�w���S���4���
�!����B��#�lx��
o�k �Pņ��+�������I#i�Śq|�����q��us�9u�ml?�x�];��{�b�c#��,v?E��l�o��N��S]�8 �_��rL�%�o-(��_\x�͖�-(��c�{�R��8y�PV��g)������	�.!�kF:�4���@��]]�3C;���P��(Vt4~ �K������̦ݤU��~���e�N����d&u�V��������r�r�Wco��4O����)A�v��n�,����л�H�BX�dkC
�*��D�o���:s8f�2��Bɦ�lr*M�����^\DR-��u�9���4KhK7�����d��hI�����yf��;����q�s�M��0�B]%������;����4%;�Z��	eH������F���nӳ��K�4�3�=s4P����O僀�^s+�4b�T%IW��\�LP�j��v�H�ow�W�����1mk̒����d��v@q`���9i�ׄ��Y����g\��{4���I6h����'ئ�D�+u��&�ӗ�V�)�2�K%���Gu�᏾��=g�&�3�.�@\����éa;��iF�[�	z��:�a�Iգ�{L�PW�RȰ�x΀� ���Lź���G�������vQ�%WR�+����S��~�w�!��_�
�5�*A&�*Ab�Xha�ON%^ji^6X�ރd���f��׫[��z�L�~cd��������2�f�
��D=T3��U�Em�Jew��)�\S"+��O�Fi�e�,������O3�P�6g���-�iR�y Q3�4��ئ0? ����(5W2�$Nԯ�?1�LM�Š��q"m�8�`S�E���\���-9�X>Z��uH�;�R_��7
� 0`lC�7O���k�����Ji�#���ꉹJ����~:�ú������g$�3��2��f��h\�����9���6�y
!�� �����/��%ML�E��R�q���kB��橧�đA�8~��N*�S�(�����k�x�G���e3�5�����t 4�Z�o�1�Ca�:��r�LL�k������ך���x�o3x(�>6�n{3%��N�a>(��e��hSL��{�7��I��0�;7	@+bJ:W�)g5���3��������1��9���[i\XVT]���-�	�L'ua砈c�@��5�:��'?O8}�0���^:A��	Cg�=�M���S�m���v��C+�2��Y����#z�O�8$÷*#�=DTdK{^�*��I���������a�6����j�0�����S8vr��T����]mͳ�^0�׏�`խǍ��W|�O�rQ9f�wa_�uQk���Ƥ(�&���w��j��_Lh��B+�L����X���զP>�:�^oy���Va ��+�O�"l(`�����y�y��k)�3z��h��҅�I��9Jּi�.�����慼��>"E�;��j��5��y��ϡ�_O�T���䌵��s!:�!c�X�X����zi>pp���,��8��n1��R���� ��ʕ�U/+ary�ZBg+ؔK����n�3P�J~mo0|��`�)S����e�d���-Y�Or���<�~��x��"W��v%�R��D_�{H���	t�YP<~�UFvymDӆJ�Ϛh�mS6G��4�d�[���L�A�"s�M#�&Tt㎢XgU&g@��������a.�0a��U��}��T��}�V�2Xc2�ׁ�d�S=U�|ً�a�qm�3n��{�+�orY4X��"ٖ�$�`~B�8�vSf��~��$KDkn��Ϯ���g�¾� �(^��,J��1!Fn�{����)���������X�ʥ#n�'sm�����Ji9�2=���]Q*	CKH�f��fv��X'�1 !V�E�>{�J����ދ8î+�����i�e��,8��	o�����A�|j]�����E�q��g��I�{���H���3�9�YA`�ѾŇ�}�N)������G�Rz8	���������L���*2��:8U���NI��D��� �S�on� � �d�&�[�p�|��h�̢\5\��G����C�?,C(�uU_�}��ؓ��z�dMՅ~��ּ�X��Ӡ%��`wp/<�Y�����-��1ua�4�4`~�r�imMN��3aq-��0����X�V�.+z�ma��T�O1k�kQ)�}}p�T��QD�%��n~"�56�r"$�����o�ʠ�^[�K˟R�~��v*����}�N�}V�&Ƿ�o�&P$"V���ܛ��Yze�_d������>U�I��� ר�P����`������e��䴨;"D:�K���%�xz�����/��N��Cn)N48;�3���;��
���믾6�Z�����F�����NY���i�yz�堿ܧ��oǻ�W+�$d�*�s?W���ͣ?�ola\H���*C�k�L�d|�|��Q:�iN��t5�{����O�gh�F��Y�l!�	�q��^�e.=�h��,��
>}v��QF-�t�����Sp�}lxE�uE%�2ӎ��Y�����/q��_���`&a�Իۯ�>^d�3M~��jQ�,��@�вK�����8�Ň���L.륖|P$��1�V���s�YM|�ő;��IV�pO��L �U�	�c�Er�o�Q�g�����ǪV�a�H�J D	l4�-������*7p���2R����_��+�z��fD�5��+0��c��=�T���jO���6`ґ�k�w�������D��4���gg�,�N��3��!:��3b�$�u��� sg!��'@Ѿ��
�� 0ۥ�X�t<�<�z����m@⃶Uq0��R�-x��J5���:��nG5�n(YA�s��h��s�"��Ӄs2l���ܪD��s�#�H�7JҮ}	���G��S�n"H%Ҽ��q�gt�-AG$Rǯc�8qݺ��{����mi�·�f�Lv���N��8�p�(�g�yLz�#HQ�E��\����K����Ko7i����f$�oҮ����s�U�S�:�Ĺ�ǅ��κGa���S�q"�k����{�d���tTt�)���O N�&w�SDm^��h�D�z %����M4�RSÇެ8ڑ�s�:s�@y�q��~�G�>D������L�9uoȗ֞��VU�!�]�H	��;���@�E9�lL2ʧxṫ�S����B3op���~m�(��o&��S=mM��^8�qTm	4�z������p����F\;>Y�M�bp�Ю�4�����wr�]n���1��#�����/=V�Z'y�hl	#,�P���/�ǉ�J���Uku��A�ys�m~��߯"~�T�Q�,�a��Z�A_�*�;�8��CC��(�RS�,/]���;+�ߍL*�x
y�A���@+���)�K�HЄƒ��/v��Z�:n�2�Ό����)4sP<�N�琡�-��b�y��v�Vj��*j\��sӞ�����
p���N[�hLA�zL����|��3ہ
B׀�L���v�ܐ���ݙP��"f�.�mzJ^m��M����~r�]QႰp��bQ��[�'��* ��b� ������B����"����v�Ί:��Ծ�	�R�b�ԁ�N��P�|�VU�d�$>�TH�n3�X� [�?����؁�����-z,�W�X(e=�T� ?�W5Ţ
���B���.���D�
�p\S�z�i�Av?���Kn��|�)A#Q��49u�Ԁ�ir'&\��D*X��˝�jݗ'ҏ|3V�CMe͏�%9<K�e9��N��a������o��0$��_��H���D������'ZI��Vr�w�0HCT�uן<TU}!�l�d*yr��m�O�|]�W�o�d�Y)��6��un\[��4	����)T�F|���ze�uJ��~uZ��)r���rW2�i������\*b���a:O���X�l�/O�cYpe���Ƒ<�7{�q�\
Q�$|*|���DuB�Dj��t��'�M��_2J�9�C�2}x�!���͓���E���x������c�4!�OU�eu~2���ec�{�����/�O���K�E:yϺ�d�,�̇x�o�l�Ľ�-�#���<�+�mH�N�.F�k�}M�d�=�K�)t���F]�u��g�Y+@��&J�+ñ�P�KC|��$�S�n�Ʀ	�b�/�ֈ��iE��b5���ՋG�ٍmH/u��y�H��d�W`�8E+n���ݗ��	��"� ����V�>iOg;���<���=��j>�%[��]E��c�w��#R�(�]Te���C�%�o����� E�M��VD�ƫ(������T�ƀQ�Ҁ��%��?-���߹��Qp����z���T��<3۬�J�
��?I;c���&~w�g�,6�	�@Ѽ0���H�S����~��w�y`,o��V	�gc�͟�^Xne�Q���R&C�4�B�RȲ/����������]+�Ȟ{o�Wl`Skz�$���z1u���<����s��@�30x�WV�j�W�g��U��;��\F;\"'��`����P�[��㷯PO�5��@������ 곃�&�B��Є{@'�Du���)���	R����������Nl���%w������8�Zo���O:��
�ӵg�$5�^@���;�G�m0er�qYj�y����:�P���*س�������FR��:�9�#�+j�3<i�ؼ�/�7���Ć~���{^�� U��d�Lÿ)~Q�(J	v!,~�V-��V�c���e�#zd X�{�{?di� �\A��se	lS���������=l�&v��@��Jkv��%7�[�DG`�9_�/��V=�ޝ�x���՗�F!��)F?1U�-4�Q�
��c�A�1�4���;�@��0��(��Che!�G��`z�,b���s��~����}���*�n���|�3T�o��?�r  ;��Ց�խ!q��<y�(��&/p�[�*Z�ۻEٸ �i���0���w?�1J�t�7��7*�����}�2r�i]V'�W�(1rA#h�:���`������:��{I{-�i�ΒF@���+�e	̬���/������j/�v�ql�0E�~K�d�U? *�$�Z�w�9�@�v?��;�wr����&����d4�B�[�hP{d�I�5��\�Fg*v4�W���X�e�6�
c�n�w5�t�I� �:�_����>n3��qV���\�Ƕ)������D
g/IC�[���(w�{�j�x�綾�T!c���X����3U��ֆ�V]�E�:��3$������0������?΃fB����HT��(M��_�rR		�gZ��Abu㋍�y�	�}�ND�5��t��5��n������쮓�����u��3��*d����ޓ�+RjB�Y�y�X��M3h*�� ��ѯ�ư��@���$�jp")�C톩�t8��Z3]O*H���ki!�߫��x�z����y��1�i�p��&�+��Znt���㎥��1��X,@��5x�j�릻h� <Ա���=��x�_Î<�j�H,�=\��y��_����s�> ��K0�
�#���Z�E�r��h1��t%�Y;�������K�p߉V�,��~yn�:b)�c�<�x��ͩ?�̧~=�W� �R��*��T�pc�#�I�C��M��y6��P�MH����%���`}n�nЪV��RR�CN�r�1�k>��E�xGB�K�ӵ��iR�A�Y>԰��UsLs��[��U	4�k5�#����d1+��������6AY�d�[~���6Ȇ����ab�U��Nx=�z/�nG�f�2-	�	�l��09�`���(��Q��e����Z� z���I��ߞ`��}���b5��eX�Ȥ������'{ڋ�8�k�-(�\�$�>��`/��y�^�Z�.\�덊�)+�$�	6+�5/!��|t��%��D,"=|#3����X�a}��ɗ��|���^?�^�u�S�"v���i@�������5%�X���[̹	G�~�N�m��.w�����M+iB��Y�.Q��r8���]7�5D��w3��ր��	�"M�����w�>=���Q̾�짹ov�B����*?���~��/�$)�6rm��m2��V!��O�`��)�r@�_3f1��}ڹ� 4�@�j�`F�.��X��S��RJ�j7�L�|�Y�����n��>���� ��4��o�v0솽θ�FY��y,R�*��T��[�MV�~�h`�Mr��h���x����S��s%�^�V͊Z�T^�d�q!%^����,zd��
�5�b���9'zI�>	)'���~z�>Ӗ�"$'GĢ��)g5z��o}���﹏6o���~R2��[� ����>B$�3�V��]���� �=�k�e`~�D+����k���G?z���q�7H�Bb��1%63TY���"ا%$-�H5���q����7�c���a=�:(J��u�E1��R����k������<P��~D�����v�����7F�f�~�u�.`�N#17ɵ��EQ!
'����0K��C[�;'�	��z���-R�c5��ڕ�j�0�e;�ZK�CĪ����j����HԤG�
3���R�G�~�k�,����>�2D��o��T����ho���$.��m6"�|�I�v;�,54�ˬ;����o� 6�:��+!4�]Mo�y���]�8kR E{�X��:.õ��ߺii����%��QuWo��&�ГbcX���,e�Ι	��r,SP����N̴�����U\��K��y3�S�T
֏�\�4}�϶�P.zE^>��C=�0m�O͞抵�%�E�Y���� zE,�$ŏ��7�����,�P^�����#�J+�T������F�,ݩ0������C�TԔ�RD�'�tY�o��"a~"B,'�w��}�� ��v��9�ͼ�a��?�8G��9�nOx��Wn^��~"�#����� 
U~qGU��Y�XH��+o�� ]r�o~��F��_��.Q)2�F��_]Y�CuQFf~v�B@R-<6,���8K�dP8x�p�����Ő�KoNk��5�6�5*ڻ��K�R�l�xr�@M��`����"䓫M�
M'� FJ��wd[MRtq�UB�h���b��n=�$�#��8��ߒ��c6���?������h0C�v��oH��ەv����{�?��k�l����;�eU!e/V[Y�?Dj�
�k��Ǭ�� �!�b��r��}��X�-\
�M驝V��7^��62��ϚkyiX�`����r�"���K�OP��$��:����w�EOi����QBN������0��`nո/C���_�X��)�ֿ*��v(�GG D������7'�;����:�+W(a�l�@2�~�}����a�~7�fb{S�.��eD�����6��_�����_�2N�B�3�Ƚ�h�K� $��H�4����ǁ�gC⫵X����r����ޗF�`�8���5�����R@ �޽~�;���R�ydrhX�ŚE2l �����2�F.�������"���B��#J�+H!M��݇� $��bg�V4����8"�/�ǂ4?b3g%W���&_�M�R��.��1���k�� "���'L湫6��O�>t��bL��"�%m��1��qs<����ŉ�H.y	�N{<�����o�h Dd��?-�����`��\�g���gV���vP̝�e��X�_HO$e���v��3�ӱ��k@�/�L�dWΨ�j�	��ێ�ڤ�;��ȟ��+���9� ��q/S�1"Y%�a:�-K�j�2��a>��#eq��i��I�9�]�U��3�msy	�X��,l�M��EB�����ݢjBkG��'@}gLyV���$So�梏�#[o˯6��:��p���� �Q����g��Ӝ��{���( ���j {`X�U��:X��^��^��:
ސ,A%���r�vU@	�L	�+*��j�����!�&;K+�.!7�p�9�\����HN�-�������u"P�PUfKaT������W�	����+%l@��~����tL�|B����1As���q��@�0"2M�&\YOa���)�!������fuX܆\��&��,R���\9��hs�t%	~���hec��	#gk2�I��Ƕg��O� �
��Q䪤#�+4� 8��E,���X$:����p����L��^�C@�q	m�B��%�&o} �cx�㳐�` ���{"cj9��2a}и���c1&�h��=Hy{5Q��4P�����{Q�x�l�>�nQ�����e��H4�{(�Є��Y�#Q6ޙM�6�0�cKZ�)5��:�)�p�����D�_����8�(��܀�[m:+��#MU�8sP��}b��Q%|��8e��4\����L<~�d�K���-Չ�'x�+3o�ė��}�+Gh��e�(:H2��16��ܳ�r�ҫ���6�zm�T�L�g�Ej;�<#��eW�5����[v]���,@��_���>Dڰ���G<"�8�	��O$��%���j���/9�cʼ�.C�V��wfΈe��@��Z�q�7���K�PZdj�i�?,`��4S[�;[�)K�W��sJ��"9�i6eI4g��UD\��qHV������c_�50�����>޲Y\���C8�J��ne���Ǎ��������s���I`a{5� 0Q�
58�y�X�F[�c��W���-������/<&�����*�ʟ���<�-)m����o6,RH]ip�� Ty�����>F}ؙ��Kɣ�	}�)UK������f|)�'�8F�9� �^���jBi�@��S;�$�J�dx��<�Bb�Q�b�+.�]��٩�'����SG���z��H����ΰv%w}�k�fl��'?p7N���c���:��,�г-�a2+Hv8�0?�3)("����&6_�~��R�CT�"9�OF�Xh�G!?p�I���KB�J�	�Z�&�$���'+�ړ]_��U
�Tmg`c\k��5�i���QQV)%�����Iam�~)^DB����+03��W����5�+:��/���)?�8#nȺK*��[>����
�E���R��9v��U�2��Uo%pCs`��Z2ۻ�L�谒�ٍ���t@�c����l��q9΃��/�k+�U���됴RU�ݻ�Wj�Mq1H��u��`&�"��e@�� �*�;�W�oPu2�N�}|�pW4��)N1kj������M'Z*]
.8q��x���q�R�����R�Ҏ�q��0a<��ҏ��	D�`�?��A��x�73�������,���m�Ә*�9a��ν
�R>�u.|A���l�%.$���O��X&5�# *�I1�Kc��]aQm�u�*�dԆ"1�~�*L�ͯd���ʌ���5��V�>j�D��P�C2꠫D ӯ�r��ʾ��z��ц%6��,Z/NZn�I`�DL��j˵��q������w�jt�g�`�}��br�X�)%����ʢ&Ӱ��La��s��X�;2$7��T�,��?~�9��l[z��ױ̮U���0w1�5X��a��>�qL�]�]��|�=˔bǒ���K�P�
	֞DYu%B��P.y�C�D�D����S�r\y�T�שx����v�|
�J
<��m��6峘�V3�*`w4/!{DL)�.�t_�ܵ�@���K��K�q#��=�f��@�}���FǤr${�>�n�"ց_&�p�)�@&�d�V��=T6�`�]F e����]�6���n4K�Q���SoB�A��v���I��؆aV�c��.q0^�K�Ԅ7�Q���i�"�f�ݔ.�~ӏ�-�
r]�	��ҍ�d�11ԉ�=M�=��ϲy)K�Z�C�t�wɡn+��m���+Z�t��po��&�>i8���Ga�1y��dw����]���\��N$+ù�Qќ�E�3R ���M�G(����.$�����" q�yH�,$<d�+9O6��z[	8���"����ݓu�X/랻��d~�$��Y�׫�H�s��`fC����0�.m�q&"���u=�$,e��������z��G:,v�H�]5b�����JR�R�v�,'A뽠|*K���E��9�zNvU���v1c�-���,Y]7�*�ݣ�c5���������M����uKu0�7r���,QY�#Q��11���/"1y�*�Ͷ�~�-fc��)0t�62 t��������eǤ&���:~��f!*:�Hh�[���6�p��{,����~�qX��@B��!&x��z ;)l>�*��[0!"s�>Q	3�u����m)��c��I�r>x���N]�c��v�^M詚��n��@��k�	��V�騇�a/���y����MiR�8���O��	���yÆ� �t{'�x��P����`/D���2�8if�g;�)1����U���~������n�[Y"0�Z$ǅ��.��EK�ĕ�BGn���k~�V��M#]����h.?��ǒ��g�z��>}����;�e<&�t�"�ד��J[m�"�*�Ϡb�\��+�|"�v��i	����*\����칫H��~2���R���@o�UJȀ�������E���Y��RQ�od���:�ɥ��Z�	�>ʠz�yiD�#A�p_�O��"�!�_�V|O]��@�s�����k:�Y�O����n6OLB���ɋ�5'7��Rٯʃ
�����"��Ϡ���Q.n�[i�>.�ek���:v��.�<"i�O�>F�ٓ>��3�V�`�kP��e5+5�vSl[�ɢ�dC�'*����,