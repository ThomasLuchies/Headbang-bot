��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k����W�z�N��VXi^�p���d�����ҋ�����6�8' G��y]A����jܦZ�����$���LB���Twj��J$QF�F�4�4s���9�	K�Ƣ,M[5���0����&�d��i���j��֨y߰YX���ҳD����@z�t���--�����k��h��y2��/�
�j9�1��Z�P=a.���R�.�U,:�e��eƻ��]UD�D���0;�/�_m��4WӇ�DK�#6Y����/@?u�3�p����rb&
U:���( v.�]����gY,W�`R��ĉ�Pה��;�l&m:�����/�h霊��1�g�9q�����A�B*pY�B��G�$Fuj֢�0�l*�1le>d(�(�(G\����T1��K����m$e��s�z�t���BL}x�����J�U����-�\*�<�c������̷���B��u�����@y d�>�il������[;y�77������ ��>�I�;$�T�-�k�\U�?B��Uuv^ֺ+,�Nde���vw[�+�<�=z9�"j�����T\�=��G�>��U��|�O.�E�����g�,.���)+�W��`S:���P=�5���FA<S�Cr�x�1U�^z־V��=����8�	$�yB�eGr�X>9`~x�jX�s� �
����PP��(�G!ɺ;:�f�,�o|д5��ܷf�E9A�-߆a�NJQ���6��e�N���0��}�~A���T�U�)�g' V�p��n?
�b7��dS�����Ֆ��&)�\!C�@Bb~����=ZM�B���~cj!�[e���AOȞ�z��?�`�$�#_�.ߦP�A����
�c�bM�547��6����n.�W�=���w#��%��s'yXʿa��ۼ���g���UV��6�n{�u2�[��.i�r��� �La�\��t�}�����j]�H���B̪0�V�S>�S�j9������hߠ2���5���^/~%�\3i�Ƃ�S�g�_�
��C{��ʀ��[ë.@q�|#HtG݇=�<��?�"��H�0̛���m�@cYT�q�d�����y��<\���ޚc5:��I��@W�5�|B�����R���_0�2nS'6MS�Kl�JSL���
�����1�W�P���
��~�a�7���2CS�8'����dS��݊�^�-"�m��I+A,������1SF{�	q"�%��=�h�����f�#F���U�_;��[a1wxB��y�ݶ���p$᲎As��bF:$�WO��5Kʂ�Z\��Lo���դ�W_�-��n|�PFe"" F�P��pv֙�A�=�;M." pԀ96��)�7k*������^d�)���V�D�g��޶1��j~-S�j:Tu�NJ�eI仔l;^G]?oW7WZ,��|׷?�Qi6�=��j4� ���k�}��|P���-�u���$�CU�	iAE�F?��婻i����2��{e<�C��/l�����#�M*�O5�4���`�� @�����*�f���v�b4��Qk�!��  a��9�i<���{ RdR%`���e�6��2%�a�$�㔩�?�!��8��� S�Q��F�buo�%��Ng��1x�L����{P��R�sĶ�װh����!�>4ɓ����q�G��iY�' |)�9��>bC5O�#4w�];i�ۣ���7T���g�ȫ��t����Q�KJY�M�N�I�3�+���(��U��,���0P8I�t��j\�>ţ��;��-OI,/����+_E+���ۈ�b��_�1.5�%zh�A�oh��=�>-(�Vt*_����5Ĺ��
��"}/!�|��Nx�`�fݫ���q�	E�vg4n���0�#�6���[-#�[!]����A��~�y)������ܜ܈9���(��'[�B�>,���� S/$^7�k��"Tva��~��ȧ�FV��2�[nTO .���"]�����!���)/�N~e!��ʨ�=��tD�պ�����{�D�x)*����X�6A<�A�D���@�4���1�����@�����>e��Lo�U�u���	�{��g���G%�ğ�n�M�y-ǀ ����/ÓFt����*�A�w���ɺ�����(B,��v�e����%L�Y�Ի�)��lh+z,�p$�H�g�f�����u�ǅ�L��)�Dx��?�O@ݢG�+#�1�Ս��˅t=�H^�$]�]�ؽahbP0��Q�����tkex)C���vGFk��QCǹ�J����6�!~s��0���s�!�	X�Z���d:P�x�,gZ="��OL��'@��mfn�`1,���.��HTS 4�K�95+2Þ-���ܯP���*97(�-��R#.�J��5Dnd�R9H���7_�@���=/T�u��]�h'|��C���날&���p�~sǃ&R��o�Drך�ֲ���0��,U�����ЫT�9���%�@8qE���LN$���aRy�(���AM��oGd���P;P�]�پt�T5Cˠ�ǘ��˿�)0�OHZY�^��Ё#�H�.r�}P�'�ᰢ�>���.W��vɰ�q������@H���=/����B�#(��&�����E��0l7�'����	0f=�� ɀ}|@�i�-�ï�7kd�{4���R5BZ�s}(rN2A��"����Q`�D������h� �OCҝ#�M�|�5��:�Z���G�4��4$�����g]��p��Ъ���6�,�6����||�~������.�P� �&��a�8C���T���u�|�Cb��gI�$��C#�z���sVp����P�#΁:���E���q�jn�׏|~��7޲��H`ݙ.1�H��^��"Uc���漃>U��=*6��=��o;�7)�Ł���a�*��[]S��2�`�>� Ԉh�B��к'~!?G����~�)��5-�T`ϋ}1F�x^\�.l��n������u��Y�}X6'�÷�F�1�G������SjsG�c�^�I�~i�[�u���2GE=׏���I 0�G��z�S�#�:3t��]��^���L�#rP��[F]�<�.�tGi*�4&�B�k�π���W�#!�c�>�M�,��]���?�8`��^I�#�\0�������}'��O�mˮ鉺i�����]l��4��.v�����Wh���,,bW�#��7G�%y,R`P^kݗ�C�Cf:��*F��j�_�w�PBf��ʜ��Հ�X!����g�'k��L��C I5�|�ʘ�YW\Yɂ�X���ͻ�Q��!���|����A����!��'�J��� �#�8�Xd8A�^"#Ǟ44\T��c��}�Ί
����t�sw�E�C�q��;D��� ���g(���q�O��̧)�� 
����lIm��M�액$d/ �v�M����a�:�R��߅�FS
�QB�]Q/��|H���A������	)�A�V~wɽ��n�B�m���?���a�Oylò�0w0)��x��ǿ66��bm~\�c�1l���zٯ���,/M[3޻�*n^�Zk!P:��mS,?��h�Fx�Ҡ9�2��Ѧb��j��y���Ջz���J���Qr�׆��{�l��'	�7XM�v�0X�kf���AF}돎0��u�d��\����Os�V��n�����W��TN��M)0l^��Z��aƣK�a���v��}D���D���= �#S�t�Z�ڀ��/��c�WҞ��w��">[H�)��N����R�Ww3�h�mOo�S�!��� `���B��P���Dn�Hȡ���ihd3�NuC��$�LS��hD���X�*RE�,�C2�+k�2������ʋw��h~��ϥ��&��n�ϧ���j���I��ٜ���<��ا�V�{�yS� �pJ�TLa��c��g�,����'���s�H}�(�!�&�B�_q�u>,���$��
I�%[�~���bpd��T�-�q��s���I����3E?�ǟ}wرȢ�#�0�"&�����UU�q)���B�D�.�H�,�j��$�u�?J67�P���m6E���G	ԅ��&	}5�*_�-�����}�`��@_�-���j*虨�"jI�����2R�O�mǉ܃��bg8Dm�t;Ш��J���o�A���?�+���E�Y�>�3o�����Q������]k��1Ӹ��Т�rʏ�._�y\�JL��*���ځU�RJ�ծO��v6C�s^"+��ΒU)ؓl������)7�q	Dg��i�z��=x�y������02 ���)��.��� ��xzT=�q�ɚB��#  �����WZx[�8�Rp�^C�%��>̓r-ӟ�3���$��O�R�ۛ�as�?:�Â���^P��k�Yf�A�M�=$�6��<���3���j�jġ�i�Ѓ�s@Z�|j���A+�.�k��8�I��Cw��B§./H%�@o̘�..�����]� �}�(���~��:�Z�!D��F�DC#��y���9�#��I�!SC���� ��	��f��ܜoSVI�x�No�h�ă��m N ��_� 3���iE�?q1t�=?��4��d��+k,�;a��s8#+���6`apXȬn�����0�1�DXجaLy�^��o����6x?#0���$How�W�_��T��א�;cDEȧ�-��>���R}�������2�X�d	��-��c	٠>}��-�m�	��BL�@e�i�$���i��d�E�/ ;�q���(��VAd�v��EE��N�^dg�s�.V|��*��_�ٌ���޼t��a����G��{**� X�q��_�dQ�9�����mp�Ի��i0#U�ْR�M�q��RjE]}�-��'n��Kq�km�m�R���]�h�tZ�y�|�e��l>e���.���b�yg��A�T\h����]�Y����lDp�ʼ}�mI���`��S��F_-ĩ0����Fm ����q���gN�wF����a�΂��͓�V��>@XR,��_�?�	+ۭM�~�8��}bWx9�@u{��h'ߺ�9�x}M�ؒ�|qV��r�L3̫Ƶ[v6�L�-z�8�l�:NRS=`�%)?���׈��Jm��z�]T�"`!�����x�&�����=]���岑�F�����hK@�����4��^ {p��l�M�I��[��_���(��}oRRE��٬��47��*<��oe)dhp�C�k8t���l�p�7!��B#�C�����K?>�!�Z��_��z��u˳?����
�U��A�D�!Ç�����H}@��=T�˛��hV�8�G5��SH��=Q�+��#�L��;aP�
���	�Gr�,�dQ��3.0_2������@ ����e:�fk�.	F�a��֩E�XL�[[�M?���7�#t�A�S3�p��7�ci�����]��py�2`N��ίS��A&ـ��5��W�|��jU �"\�JE���R��1mF��D� ��*�l�蒃�Q(uٛy�ό�7��I��sqvn��ԧ]%g�;��QfeΈ�2V1�������mT�;\"�n�9׸�E��t҆IS#��Z�L�`J�����hڿ~șG���N�s8�����o�ϚU�{
�/I�E��Qr����_!����K��UV=@Sh�iއ�|�
����}!,���["��<U�m���6����������AkBk��������;�0�����ո6,)	�ǫ4��R�ȏFrCj���i'33�Z���᧖~0M���}:uh�{�DNH �5�3Ɩn.u$�#��O���$,m���S좏������3�5c����b�ǋ9/�N�o ^,�QW\��^t����m�����	�_(��Te"3l�kQ���+�e��k*�,��ix��SS����pT�"�J��]�sg�W���`��i�cRF��Fzv�m�+SLA
U�9N���r0�^k�{��f׽V�z=a��-�+��c�����_�IzQ�\�x����)���P��xǿ��޶���!��v	7���D���Ug�yeK@��g�P�?���~����WJB���q�y�)�Ib�`OMn`�R_�	퓸�ǎRw�^��0F���֫ =�&�A1�8���n8_����ځ�����o��IE?mR�jr62��L�����������K�UnMUs�*0I�_I��U�Xc���^	�׶��2v]o�P{�9	��ː33���ؕ�:��~1����+�(~O��)�ym�X�*�\5N�>s�]_�#Ib�6LJ!&f����O�0�w������ͧ	[��e	�k^wHJ�-o�P�6���A��c"��(h��vpW��
)^�� '	���({���5�g��LI^���ur\fLV�c�C��F�����w�ex��;�A<���Z �A�q�c,���Ò�,c;�����uN��+GRܪ=کA�7Z��
�f���k��.?�h~���h@�(n����*�\��p�{��M`1����	�2Ӝ�OH����!�[Ɣ�V������ONxIe��ƓY�\�j-� ��މ��A�"����A�ƫF�j0�9#����O,Q���	���rko9���S�L�a���_r��,T��^C�y0"��d��?ڕ\�����Ъ/��&߉�����*���0⸔8��e�,���we8�\�C_EL8�F=���F��B����9��9�&�탴m�f�L@������h�����ۧ�o�	D]�=��h�-6��6*�H#��"\�~D�R������W�J`��E
�'X��[g�������X���%8п�*�Kf��<^�D3x����+m�i�)��җ=mE�J͔�'��$-��o�)Fiݫg/��U�n}�s�T/�]�h̨v�+,g�Z>'�5ݲ����0�c6K�!Kh����̃6�r�=yƈ�������w�59��6b��5�@�n����)�����O�:�3����FI+tįp����+t�R�N�*�V��75�]HFp���xp\�N9s)�&�b�E�-Q;�R���~%X�sN�L���h���:L5,�S	��S�i�.���� PУ��#N`�^֬��ܭ��6>�f?Q��
�md8m|�<��`�b��!�/���\߀.+Diw��K_������]Nɛt�������w���5A;Q�I!r#E��΁%��+n��~���<<+��'S���g<1��j�e)"��p����9��CeMh?������1�6I(d-n?�S��`#>�6��[��x�;^�焽4f͹�d|�D�8�|z��N8�@L&�	9�ֲ�39K&By�R\���u�b�Ky$�,Z;Ѯémr�� �b.�X��`��_����+wo��<ti	�.3���ϓ�o
q|�����y,0��;:A����������ia;{ii��Ll�*�8k����L�"ţ�`�G\�.��Ts���:��*��/}R�\�w�� �x3
��ұJb�*K�]����Z����B�ed@���5����I��^K�F9Js�C����2��,J��'
�h{a.})u=2��o�i�����h�c����i���p��%�����*nj�ۜ�i�����T?洼���4�m�LB��g�����n�~|hv^A1v��*o�:Dw���X_~��$�"�Q�/������%�"���L�ff���C��D���O��[�c���Z�k&�R<�#�pE�SH�c\!?��U�eWӷ��ѭ�&��Tf..�))�5b�Q�Ǎ���_g6�Vk��Sᜐ��B���1��S��j�!A����IX����V���"�ė��o�����i����vv�C�w���xi��F����ρ�k�eI�!���f��
�w[�{
�Z��鷶��s˄+:��rФVO�"��(��|3 ����5�K��"� �����WSI��i�Mi�j�w�����u�Ɠ��ǄͶ�Zt�R��dE���KVs?*�P����vz����Ԧ�|��ּ�*[��b�ϯ0��u�V��E�R�h�y��g����.�7�
�v�����Oä�7;�	�AA�6p7��˵�󈞵|Y�.9)a�?�TO��OH�>�E`�����0��Ղ0�Nu�tu�/	*�/��k5JSVN��(����3�\�ᳶ-�R�&0l҇ ΃�J��gg,C:9�C#�Ƶ,�Riʃ�ޭ)�t-�]�ٖ�y��c��c>�/�?,�����x��"�aUN���%l~�
Ąn�t��ق���z��rK��oE�ʔɷAs����8�U��F�D�&���0]���$^(�����f ����:~b�ߋo�#��s��0���FC9���W���0�8S8��+�j��)􄶢�fo��>�\D������8��d��_f�-,�v�v�{��4�g?��x�ˑ�)˽^����K��\3<'�Jd�5ZE�<8u�k���Yr)nO��5�h|�-x%]���T+tK��C��9J������ǸZ(�,{.h��tG��eKN�^QL�6�\6.]*H��o���@���ਪ:K5g�@�˺k`A�B70�k��IR��"�61�q�5b���
��,#H֗����>sJ����wS&b���}Z�@R.cp��ʁ�A	j9����X(\�%8m�O����Z��4N;��S�Y��yC�i��X�����}G����k�bW)#|�%�2t �O�7k���*k�+�?UF��MtF�L�WS|�5R�nVi�AZ��;�S�����N�>l��W�;mik�v��N\�vm>+�ZB��<S�~�Z���ݫ-��F���
�����E�Q�z�S�Vnzt̃պ1���b�>����O�>�d!O�ĵ�=�2�D�J�\��H֝��*���2)&�\�trr�a���^�zZ��B�ϻm��$i�ƍ�d�MߍD�R(����4��x�8��)o������#ib�{��;�n�|sr��_�+���9��Jk���h }�!.�I��I�8Xu=�jˣ�J�Qq��5�����eYhNJ� �{�L�ň�?���!%J�X�#�-\�TgJ���}� �fr�
(��l�m)�82c_�^q�|��ǘp����X�W��&�C���&��t�je��|X�Mv4mk�0\�\�)�a8�Lg��[�4��$�5�fc+jM�,%9�w��2��rA�ZPL<ֽ����ҩ��̵�pK-c��!�O�td�i{=y�gwŎǖ�X�K�yq�.\�7��
".4C���9�q�Z�2���.k:x�������������GO���6���Yޤ�!���X�f
z�B�"_�߀�.�"pGU&��]k�@^
���m[#:8��=��B� kn�q�E�0���}�Zx�N� @}��g�a����\9��q{_�s�ͧ��v��[�;>3�X��1n��(�����Q����f�"E���M��Qo
�wt{4ݕ�~�~p
,)RX��@��_R��)�O��ׅ̾�� ,���s�s��#�[��d�)�!Q����%=��^.9� �2��B#U9���J�:ܞP[��	��HR�J5�O�\�.���J�N�ǩ���z=}���)a�s��I���m�6��!��ϗ��0������ۃn��� ](nsܿ�C�I(:)QEG�i�����1޷�;�y�PWWQ��F�_������N�O'9�s�������P ��m6�04Lئ��P/^-�
xw	��C�s���m\ld!�2�e�-�RXy���^�t���-���Q�]���9�#���Y�t��F��|6�/}Hߦ���s�+=�+�{o@A]N�A���T���Q�H�e���'��+޸n��a��Ӗ�k~�B*	�,ϠK-����6Jv�h��DV<�C�7�o�kKFx��V?f�A<2ȔO�ܘ1����thH����r9�r������.I�y��Jd�p�_xD�t�C)u��	C��L�I?9=���T��N !6K�ֿ{�������"�iC�(�M��'3e��y�#GwT��3�	8u+դ���n����%���Ҋ͇%���M�F[�9&������~N$I3|v2#p�����yb�m��O�a2����1�����NO�,/���.Dc�b�`��^��@�V2�	&�?�	5��(�n� �1�$��z�����	v"�۲��F[��N-��"�t��K�sr��A�l�ét�h��o��_N�>���.�S�<�H��ts��'l �BHE�B�N��W����Hc�"�5��9�{⡃�kҡk�����~�IU���TM7nE?>�;1����A^��k��F�M����$��;ݱ�8���m���fz�K��"�ތ�UM��^����~/� 8`l���`�듔Ɵ8���������o�N�[_j��|��L�3B��a������t�����k+"j(-�{�#�����ykt��b/|���v��	N��s���2-qcJ��m���^K*O��,?�Yp���ӊ����^̇�����	�>h����)��z��䃚�Vrg�\�uS���2�N�0�n|)���Q��o-��u\��>�qD×�C��^�5^�%>��k�ڤ*e�ۘ0�["�^� t7;I�̾��3ӟ.��=%�=�X���b6�U��a7���ׄą� wAxM<�W�&Sɨ�.(�9O?��!����gQ���CU1���j��@�cd�OݠW��Ն���6vr`H�y�θr��d����*tj���	��!����|�����P<��V0�Bm�,%P)V��Zm��W����á�̮� �H?nd�~�ex��FҀ��A=�f	x���A�=H�W)������2�smHc.���.#o"M!2J�����hV����p� VX��v�o��L��P�K_���*١z�aM��ޣ� �`�m8�������:��&b�<7�@t��m�p�޿��H�?P�un/�$R�V
�׊�[���Z�d�X�}k1g���F�&ܖEIi�V$���$GA��؄�ot0��3I)�|Q�Dj�Ɣ �en� �m鍻gҜ�2������:,=sj'���y�­��$���</�b�aTJ��W������O�,�9i���7�u�e���|LS�x������p�R�y����U��.�]�ς�iP�8���
����i��l�i�q;W���Ƞ����7�T`2��,�z�:��� ,0�vο���ِ.R@���F����������r��mó:�7VA�����w{�<����k������lB��V-�sd��G8�	���l�
�Ż����gw*�<iY�Qk��k���[	P3�Mħ�^��ч����������_9@���#�!����A�ohm%�L�Ru�8W"����.�9�P�=��׬�4�1������N�$)c�fW/j�|����z	堻���}w�ќs���˩�.^�7ik@�h���H��e�P`�����"��=��ėn��5@� ����>p���|�}��{WDG�"�FC�=B�E%�%3ee��x��D�W��fF�����)�$��Z"�����?>H�����~�}�nyZ96[(���yy	�������@���/�!
e!C�z�M��ʠ��[D�1�s�� ^�~jʬ̚9A[���F����	����d6��&5�Z��z�!N���E�Z�Јe`�b�(�)� �H����)��f�ڔ�f��7����i���V��Y��"��)g\���]ǰ��z�1V�T���zP�,kM��pC:����Ml���d|��Kc_�,9hǼ����+�D)��P�+�{�$�I)�:b��XgV��Z�+��pə`^��#6I�1��}���f�Ɯ����X�6�d�^is���?ŵ���eQ���8&v~i��7��\�)m��4�7��8G���9�V������	�h�p�F�<��+M6"�����n׼��C��z�hg��l�e�F[�V�p��ҰI���s��ejPk��A~(�E��[@�B�0�r�B
;ǅ>�PF��*^N�hx	P��f�/�g�Za3�nX-S�+%%��sqq�O��Ϫ�l`C�ȁ���KԊ�^�a�:���ÆVa�$���<�)��/��M�=��������+�=�!�q�?�f����N�&�zŲ����̙̲|���[�7����"$J��X�Hf��	��֯�ʵ��������<3o��O#�j�G�T���r����J�_����9�q/*��2�����8v������	gb>FO�g��0x�>�,5�X�⫧q�������Tb�Nкc��8�zL��X:�4�vx��;�7�C�vw~�Pm����Ӄ��we���0��W����G�r��g�w��O��5�[���
W9(�y# �=o��8h6��(����h�J�q�%;6�H>��+򊩵�I#�w�s�N�4���	O�4�Lّ�o�@�3����pz�F������K"��i4C%���I��ـdr��$��XN�ωK(��n��w�%���ް���КiU#�j��ː��٧�!@hk�%iu�?9E(�c�ӅuA�_�N�0OK�7�\�F��+8�LB&ګ��&���v�H���(CG���ET��c�(�#�fo�\���:OM�jb�,,ܛz�	�Ӻᢾ��:&�N8 �ͬ�>��/Hs���������0_��zp��\�r!�U��e��bϱ��C&~�Rl�M�9^|��6�?-��X�n����S�����X)m:���-��J%�Z�JI�b�De�������vB��F��"O�J�V#;��ًu�M�?P%�'�-��G���LZR�j"���ez�]�k,�ML>�� o�s�J��a�=)f��%r��`��V��7'&*�6��n����,5�_���-S���}�����F0�w$�{Μ��Y��Am�h��h�K˶פ�G�5۹��Y��؊�|P��G��p�s?%�]e��켈����þdHۼ%_�4���ap��gρtato���5ou���ʱ"�k�;p|p�]��<�s1c�~'_�ֺcZGi���۷Ӽu�9~a8�ڡs���SZ���!B��9Tx�	��4a�.t��Y6�=�@����.
���Ϩg���?^�S-ѡ�aњF0��
ķW'����#EM��?�/��Kw�&6��.�ǚt>~��%ʋ���kC;�Ե�j��`>������t��!Z(�Ĳ[r�P��Y�`$�r}c-�
	�G�v�� �0���Ƕ�����%i���<����یVu��#U�W����]��BL�=��N�`�'���Bl��I:����S�n"��)�Hh�<a��t��yN�v
�.�N �6銶�Wٞ���r7��
�W���Y�6�h��N���3�;�``(Vq�����x/a�q�b �*Zx�<{�!$���x��"S�%s��{6,����猌�K%i��8slKv��p6��F'[�ʼ5;&0���J��9�@ ō�^�E�����VVj����/y5�VB���~�������^�~d8��2��B�,!�G��l�'����`<���g�\� L��n�󗦎���e���a�EG����v{�F��[�����hL��x@�裺,\L0�X7[8&�m�IN=�x��v��);t�]I)n���Y/bʙiU򪏳pt��ts�f�_����JZO�Gʨ�6I���E�FU���K/��@��"�,3�K�L���"~k�Jŉ�ud��3e���.;���a7:Hg�O�8Ǌ��M&/�F�zZ�+��F_�A���-���9U±���#+%#e�eXs�pe�c�`G��F���*oҋ��jaT�e�E1,f��?J^��x�����с@��cTŦ@�l���c'�s�V1�qv��w�P��αO��G��[w ���T�T?C3��2���<��T���)Wt��`:��z�����H_��R��ӭXUQ�09l2dw})	�Q���Ho�N3��̇"�7n���R����ޠ��(an`�T2C=�>�{Cż�g��9E����4R�I�[�D���r$�ũ�v���Ā.�x��0�xNU�	�C���ZEC����`㷐#1��U�o��o����������mL=�UH�z�]��N����[7o��d�kd�xu¹	"�Z�f�\~���xV�\G�L��B� a�����! ��62��svo�(r���i��-y�3^��h�@�*0�kRC��~���5��}��(f�o,��'`��}��2XJ=0������y�0t������p�N�7���"d�*�O7��#O���/j��L9�ar3�2b���Y䖻�t�nε��O��&��w����{x��E3^�K��?u)�?z����z��p(C�o��O��%ZV���6�A� ���|�0�]��Q���
���I8�a���~L�5�}��t�����ҟ�ډ@n��P[J%�ॖ_��{�.��{�`�H|�2���%SZ6E0U�_5#�V|p��Bs��%�_����L���zϸ@�}f�}(�h�.�J�$��U���M�S��ǻG��N�����I8G��/��\�	Z=��\k��R�a=����H��+���	�S���*�6@�K�XGnY^+68�γ7��1J�@ Oׇ��X�Uѽ]��`�GBn\ 09$���z�NX�gnL%��xm㹜�kP��p��e!��ٕ���d��H���^���vͬ��fj)�R~�j����F�>�+:~D[����-��ϡ�,ژ��'�N�PLL'ҍ��E�W�A>����7�ʩe
i-<����g� �\ž�O��,��¦
H���M/�7��+�d���f�[��Mi�^��h����y�H��A�Ϛ�Qѝ�w�B~�'A*A�q[:���2����*&t�2������X;Y�rW���ҝ�ГM��@�œ=��'�?I�3r0���B��
4�R����kE�s������k����x��8�/��� |Q�s<�*�m����ة�Z,�J�0x���)e�������H$��]:��M�6�r��NՂ���9��B��M�,���.cx��Rg�u��&�����B�\|�Qs>�!!�&��g�1�C?�)Ԧ�]Zd��q= �\B�u40�9��~�=�.�{���B��zBx�S�Cv�۳um�v�:%�ӆQvgі��=�=�&��(?	}6��L0D�#��f�ԙ�JV�������L�R�ɳ�;�v���{�w e��M|��^KlN{o��ؠ;��m�cI��4�MQ'n�3��}��Q�&�	d=���=��E�a�/��.8\�B^�K� ��cC> I�݈h뤸����ҭI�����Y�C�j�B"�K��Q�gvI@�� $ܺ��{G9�w�2��NCP�0��&���hDJ�)��-����d�k(�-��s?|$�Xva��(����� �yo�cO0T�o+J��}�6+`&Y�=A������V��l�-B�#}���: =�-�1�����<����md�- �Ha<�zC��ު䌭�,�#Yhp��O'�F��g���]Ϣ$y-~ND|0g���ҟ���ñnT�;�UF-�_��%)V�T� �{�)?c�K�aLO^��&U��E�����s�1�� ytAA����F���T!�rU��Ltz$�W����H��1n>�	��A~�[T)���!�Ja7(�!�zV�ǁ�^�פ�����H��jK�N8�(��T�B�U����g@>�KO��>���Kx� �� ��,إy
�Iξ�a�����k4
�b�gfR[����Ϭ�1_S4I�`Ѻ����uą��;��� �v�NW�ü��5��)���Qo�`�V��(��Ä�55�x��J���X-���Zȃ���������M(�����`�!2#�=�|�"�_�ձ�F�����ۢ8�v! }���*š��Q�kS }7)�C��%��^3������+� lKTL&���P[=#��srO:����
<3v��!�z����u���į�u �М�#���&��BK�?`*	���h��������v#�:dڌ=[;w%��ۗ���sq*�>����,9_�6�����c)C���x���0��\�ސ��'R@������p���)�㤔�����U�����M�m�@��*&��J�y�ݺ�I0��jG��m��Z��$E�b����
�x��~̼׈4T�!O-����3(8<�X�,�qo'q�Q�w*��'�����qHM ^�cЂ�_�fq^�w�h��y���k��I��\�:g؋�x;vX�/��V�6�bV4В�Rm����M����稀["�.F>]·-w���$RBkS�(`��[��}$Goѫc�+��گ9�Q� 1S�p�H�$pn�������G��.@�?�RpN�݆�Z�� ;(�I��'m��03),����͎��O�Ǒ�G�k7���٩�3�5V�j�P�V�(
F��m��2�k����x%�@��V^<��ƹ�<R�%���+Շ(7�+���=�%)���'�7�����(����%��#e�RK���y睍���XC�f'���H;<�&b�½�g��J��ćf@����x��nVq��y@�3m گ�	�3�BZ�&���������V�z�T(��i���u�GX�������|'A�y���O�K�c��nph��:�����(D�.v��\w˔a��s$.���Z]�������Eu})�
�`��`x6�\�N�6Bd�J�x遜\��S	a�H����Kw��N�@d�ɭt�iզ��)�N}�q�����~�\-B	]V�(D{Ȗ~�ﲽ�s�/}�h'�6��kI�X_|�;��դB����&�f<Nx���	���n[I�,�R+�a�;�E�I���7�bBr��05 � `��X��GY�|Q�}��2�f��;���(LBY�Rx�������LR�%,�;ĵl��r��vyDގ0�����C.�ģG�7����x���]���¼���#*�#B)�;ۑ�w,Sw/�F����ҝХ��f]�ڍ�,�VyB���� ���I�W�����
��S,�`UC��_��2�<�ڧ��U��=���h��*�7Ur�U]��ۑ[��A��H�wlw���	����@���8O�
�f(�`��`�2N�����w�Q�(�p%�GCk�Ѱ�6�|��3Y8�� �2 Ý�q��8M�`�5ϧ5����ҏ#�HM.8�T�1+�̪�*B���8�(WRp�����j�I�=zE��b(�Ŏ�eL�r@۩@��uʲ��Q��q� Oi&�A���:�"8������T4��<{Z�!)�hB�����3��0	,\�ϸ��]�L7��A��;`��\���m�E�ZE�M������f�y�#4��}��8m�I��Ȓ��z����4(�c��;��%�ܝ<���S.�O7���F�>���^�����	����N�[�����ox�`�veN���0?CGg��#L~��4�4&���k^���K���N�H��wĸv�-����IB3�_���S^�����$�T�l���J��p�i�
P�� ޲S�&'�nB����7h�i��F䵑}��f3	�c�m �e�N��5Ѷ�| 9\�����W]�C�2a���=v�C�؉X�F�m�0 h�:�>yQ��e��0�A�+�j���5�������G�\�/Em�$����Q����K�˻1�f���Y'f1��({�|YB��(
��,�l#�N�;2��V�ȾK#%&�5�����a8���'$�����!� �˰�J��sJ��p��\j��G����P���^+�	�h$����4�C�7�6�y�k�x�57G�,<����g�8���?%�����U
�*�w���Qc32T��C�A1��!c������Z��@����!�v~�{ڟ��y����U��삔O��7VY�L���6��m�&E�
�!�%J!����m<�����*�?F��>Ĵ+���Q�4�i=����і�c�7kMT�әM�\s����`�-��AZ͐sz�i]t�An��gم f�%����Xҽю}Ƌb��Dfg�'�P��$�<3fSX(8âc��q�K�Ӧ`i��*�ԏJ����Y��@��L�*�'k��5K���uvsk�9f=�՝�rmB3�Ϙ�<#�s��tT�erBg��Q*�T�Ͻ��*{\�@v���z)�b*.~����N�|�
R'��'����) "o�`���b3z&ו;�Ρ���Q��-�r=�t���a��p�:�gH��Ѱ�����PkRI�H��l�������Ь�Ɗ�*�K�X2$�2��G�w���ܗ��*�������Ie��wJ�NZڨ!��C�X.C	�����hES����P�9ME�����f$��I>��U���z��_wݙzS�1[��53�p�}����a��y��>҂`�u�e�9��� ndu^�@�䊎�B2`yB�F�a�L�c�&�k�SH�{i&d�|�VC�C�f�{?s� X�ù�%s�è�����GYV�l��Z���Ccb�b�����D�����5�+�����#ڃ&�_�`��{�X��?
������O�l��Ç��.L�6��y_���@�n������f(�d"v�?0#$ _��9�X��"1�U=EM��+@+�~�=�R6CM�5Gl���s̈5,�|As��]��Z6���1Y��53_��ఽ�b+c��W�q�oLy�@��>��W҇���f?��k�Tz���W/�P�q(6cR���	y��kã���^�v�U@r�4=�;J�܌�Iw�g�Y�{��A���}C��yE�aJps�)kZ�{Q���$�o�E�i��Ϗ?��xT�"�I0�;l�*V�ۮ�	=��FZ�5�����!���*ˁ���K�Ϫ�V�E��y#B:ǋ�4�F�?�=W�տ-����LP�"Z�|N���~v�.&�������Z`_�qb��ֺG��X4����Q��`�	�X�ɔ̶�*��[gu���5`��q7��1N�	����2�|{�J4����$e�	�,s�q>��iy�؀>��	wкV-���!X����tpK�0�?J�Ȅv_nJ�c��	��H��K�\w|�#�/n��`���5�%�6��i�����L�-�J�&��yՖ���@��Ԏ�D���$Οm����l��V��UV����	��\Z���ؐBC9�%혶t1B���h�Z����TU��3��䞦������rU�)���	�(&�,�;�W�����{c��G���]���b�UB3q��D6O����9�f�7<����9�$�g�ꐅ"x�*:ռЪ��P�3Q-���Ǵ�X)R����Q%�E�<2*���\ᯊ^}�������xѠ�����(�fj����o'�+�7�\<O�+^��U16[ɶ��8E��{r��1�ƀN��M,ش4��4�#B���'���{0�n"�Z��ڿFN�P:'����0�[� �d0�=9@�B����Y❨V�ϓ�*��w���SgM�$���n���/"�R^�:�y	��tP�=��s�52��#Ӷ��r��實|����%?���.fI-.e^ �ŷr;�u[[f������i�A֑(�A�\z6���ũ؍Գ�o��V^j�[k��]�Z��Ԛ������'����A�-v-S0uΥJfPO��9����To�O�����Z�MC����kh�1Ebd�i�`�LZ%A��s)��˻��6��3��q�X�E25ܦ:'5���� 1��ɀ�وZ��S�7nٟ_k? Ո��f�Ջ���/�C��Mz*9�ۥ��I��RO��ci����SW�+x�N��`��k����价3Х�@YCD�O��rt�h����:@�����,F0qb���U$��B�����4�ʳ1����[Y�~�f"��te� :���HJ\�C���G���L�^*h���WY���������F���I�P`o��m�w_}��o�VT�C�B��>�	E�{<t��b9�MQ��z��=��2��+�'�b��C�d5� e�V`�z��wP� b3����H�ѡ��w�f{��5�֓L��RuV�s��|���.LCf�Rqs�;�GBo#���!�����Q�׬�0\e��xN{]�ga���Y�C�\ 	lĠ�+X���&�����@�e�c.���w�3y�?���.�����DO�����H�^��?b�.��.��`á��$ Z*	Nl���`J�����ׂj���%7j�3�F�F�����	�2c�-�-�q�yDpw����o�����|�0����k趺J�x`JހCհFaSeMxa��.x���N3!�g���pȋ�-�hS�Ɇ���a2�8�x��P��Y���D��b���#��d�MJ�8�VKm���/}�&�ܵ$�񔋂)��� Jxg���q���1���yO^�>�KN��b*�K[.�� J)���md���s&���̌G0����|��^>�Cr�j�	/��À~����,"�`̫�\з)�M�Ւ�L��~��W僿DD������v8�-��g����j����<(r��eQy�'R�I����͐"K쪿�����/Y+�$�_!�b!�9���OL/s���K�ù���Js�����E��O��Q vP�e ����T~���*�W�2~�y�Y��@	��0�.ՙZ�=��7�3h��js�I�U�-��~��<~.��c��� 6R�7c)�����f\50��j�P���i,�Ϙ��R-�N�}j��pɻa�J��r��-���Nfʘ���[Jfn�t���l,M�\ܿ�I��X��]�d���F�� %��D_X�#��_8'�Y��~h�α�<,���+�~,f���t��1ؠR/�t��n6k
��Ԫn��ս$��Z��*�<*�Y�뷺_=�787��'�&e�=�!�n'rk���O>{�ΡS����߸ciF�v���Yy�l���E8B�LT��9�f�r�b�O�!͛ʺ�N�N�j6���oL<t�70Cńv)�(b#�c�z]�O��n��b���ݙ>R����g�Y+w}��Q(�퉞�M������p�SX�nD�Ck�O��w��\�mŸ2,��aV5�,/S�(��D�$�ڹ�H��ɽ+�.����)H�2��CЈ��O����r��z��m��Gra�~,�i�m�m�P��<��R6RG"�i�|����BY��h��
�R�gJР�.rT:������� �ge�X/��ݣ��X)��T[&���6Bx*��H�l�,R�`�'���T�]�-���iV����Q���7(�:������0 ���3�oB�D3i<#�uL���yi��la��g�C7��RS��~���'Q;*�����xa_��d�m��k��r���|�6���tk+�����9���AO:�3��s��ꔳA��2���A�b�.���l�ێ�RmM��:��FCӈ���:�sQ�`�I�}��|���^>�V���t<-�g��鯲���7�r���v5r�V�q����4��])҂���_��鉵�k�^���\�^v�M
��1���Dg��yzB '2�!@�[@yHg�uJ�"�=��a:��e]Wn(��#᠐������F�{��, 2�����g0pmU���nr�E��	є��k���J��Mx�S;Q���P�M�k��.��#NFG�h�I�� 7����^>�安��[PV�_�xSB���,!x�hj;��I��bM�k��1�"x������<-Px�3�F��R��x��5���C���䴛�R?CV����st1�@-	��r�{8�e�x�x���GvBD����d����ڡ��%�`N���P=C�%*�,��0P'�c��b�E�(�LO���o!e��,?�e�D�>�m����Ŭo� �D��j%J&����)��\MW'i��R��0H��AJ�5����������#�	6Eǔ�k��t#�j�s]t��������P���߉m���5�]0k2����ulz��x��p!Ϸ��k�1�{rW�,�7g�s�aN��@���*��^�����������F^d�u)��Bi��n�4�k�X7�z{�C����b�������Ha+'�|�����n���7���鮶P#ȚA�����)�m�1����r��X������ڗ�#z��ͼ
^��N��|&�4�^��-(Y�����w�5^v��%���h\��
��D��� �����xOƒ��]�~����0��ўΦMvjnޕx~�\שY6�3I��0t�F>5���^���?�Uev�k����A):�	fr�n�ZC��X.��]�