entity servo_controller is
	port(clk: in std_logic);
end entity

architecture servo_controller_arch of servo_controller is
begin
	process(clk)
	begin
		
	end process;
end architecture;